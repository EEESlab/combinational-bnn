/* Module: data
 * Author: Manuele Rusci - manuele.rusci@unibo.it
 * Description: BNN net64 model stimulus.
 */

 module data
(
	output logic [99:0][63:0][63:0] input_o
);
assign input_o[0] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000001111111110000000000000000000,64'b0000000000000000000000000000000000000001011111100000000000000000,64'b0000000000000000000000000000000000000011111111110000000000000000,64'b0000000000000000000000000000000000000011000000000000000000000000,64'b0000000000000000000000000000000000001001111100000000000000000000,64'b0000000000000000000000000000000000001000111110000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000101100000000000000000000000000000,64'b0000000000000000000000000001111111111100000000000000000000000000,64'b0000000000000000000000000011111111111111100111000000000000000000,64'b0000000000000000000000000111111111111111111001000000000000000000,64'b0000000000000000000000001110111111111111110000000000000000000000,64'b0000000000000000000000000011111111111111111000000000000000000000,64'b0000000000000000000000000001101100000111100000000000000000000000,64'b0000000000000000000000000000110000000111000000000000000000000000,64'b0000000000000000000000000000000000111111000000000000000000000000,64'b0000000000000000000000000000000000011110000000000000000000000000,64'b0000000000000000000000000000000000001000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000001100100000000000000000000000,64'b0000000000000000000000000000000000111110000000000000000000000000,64'b0000000000000000000000000000000000111110000000000000000000000000,64'b0000000000000000000000000000000000000100000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000001000000000000000000000000,64'b0000000000000000000000000000000000001111110000000000000000000000,64'b0000000000000000000000000000000000000111110000000000000000000000,64'b0000000000000000000000000000000000100001111100000000000000000000,64'b0000000000000000000000000000000000000000111100000000000000000000,64'b0000000000000000000000000000000000000100001110000000000000000000,64'b0000000000000000000000000000000000001000111100000000000000000000,64'b0000000000000000000000000000000000000011111000000000000000000000,64'b0000000000000111111111111111110000000001110000010000001100000000,64'b0000000000000000000000000000000000000100000001101111111111110000,64'b0000000001111111111111111111111110000000000000011000000000000111,64'b0000000000000000000000001111111011110110100000000111111111111111,64'b1110000000000000110000000000000011010110100000000001111111100000,64'b0000000000000000000000000000000011010111100001011001111100000011,64'b0000000000000000000000000000000000110000100000000000011111111111,64'b0000000000000000000000000000000000001100000000011111111111111111,64'b0000000000000000000000000000000011111100000000111111111110000011,64'b0000000000000000000000000000000011111110000011110000000000010000,64'b0000000000000000000000000000000011001111111111110011111111111000,64'b0000000000000000000000000000000001111111000000000111111111111100,64'b0000000000000000000000000000000111111100111111111100001110111100,64'b0000000000000000000000000000000010000000111111111100010000011100,64'b0000000000000000000000000000111001111111001111111100000000001110,64'b0000000000001111110001100000000001111110000000000111111111111111,64'b0000000000011111000111110111111110000000000000000100001011111110,64'b0000000000011111111110001111111110000000000000011111111111111111,64'b0000000000111111111100001110000000000000000000000000111111111111};
assign input_o[1] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000011111111000000000000000,64'b0000000000000000000000000000000000000000001111111100000000000000,64'b0000000000000000000000000000000000000000000001101100000000000011,64'b0000000000000000000000000000000000000000000000000000000000000011,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000001000011111000000000011,64'b0000000000000000000000000000000000000000001100000110000000000001,64'b0000000000000000000000000000000000000000001111111000000000000001,64'b0000000000000000000000000000000000000000000011111100000000000000,64'b0000000000000000000000000000000000000000000000111000000111111100,64'b0000000000000000000000000000000000000000000000000000000111111111,64'b0000000000000000000000000000000000000000000000000000000001100000,64'b0000000000000000000000000000000000000000000000000000000000001000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000010000000,64'b0000000000000000000000000000000000000000000000000000000001111110,64'b0000000000000000000000000000000000000000000000111000011111111111,64'b0000000000000000000000000000000000000000000000000000111111110000,64'b0000000000000000000000000000000000000000100001111111100000000000,64'b1111100000000000000000000110000000000000011111111111000000000000,64'b1110110000000000000000000000000000001000100111000000000000000000,64'b0000000000000000000000000000000011111111110000000000000000000000,64'b1111100000000000000000000111000111111111111000000000000000000000,64'b0000000000000000000100000000000111000111111100000000000000000000,64'b0000000000000000000110001111110011111111111100000000000000000000,64'b0000000000000000000011000111010001111111111100000000000000000000,64'b0000000000000000100011000000010000111011011100000000000000000000,64'b0000000000000111100110000000010010001110011000000000000000000000,64'b0000000000000100100110000000000111000000011100000000000000000000,64'b0111110001000011100000000000000111000111101100000000000000000000,64'b1111000101000000100000000000000111100111110000000000000000000000,64'b1000000011000000100000000000000111101111110000000000000000000000,64'b1001000011001000100000000000000011111111000000000000000000000000,64'b1001001011001000100000000000000111111111000000000000000000000000,64'b1001101011001110000000000000000111111111000000000000000000000000,64'b1001011011011100000000000000000111101110000000000000000000000000,64'b1000001000111000000000000000000111111100000000000000000000000000,64'b0000000100000000000000000000000111011000000000000000000000000000,64'b0000000000000000000000000000000111111000000000000000000000000000,64'b0000000001000000000000000000001110110000000000000000000000000000,64'b0000001000000000000000000000001111010000000000000000000000000000,64'b0000001000000000000000000000011111000000000000000000000000000000,64'b0000000000000000000000000000011111000000000000000000000000000001,64'b0000000000000000000000000000011111000000000000000000000000000011,64'b0000000000000000000000000000011011000000000000000000000000111111,64'b0000000000000000000000000000000111000000000000000000000001111111,64'b1000000000000000000000000000110011000000000000000000011111101111,64'b0000000000000000000000000000000000000000000000000111111100000111,64'b0000000000000000000000000000000000000000000000011111110000000000,64'b0000000000000000000000000000000000000000000000111110000000000000,64'b0000000000000000000000000000000000000000000001111000011110000000,64'b0000000000000000000000000000000000000000011111100010010000000000,64'b0000000000000000000000000000000000000001111000111100000000000000,64'b0000000000000000000000000000000000000000000000100000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000111110000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000111110000000000000000000000000000000000000,64'b0000000000000000000011111100001000000000000000000000000000000000,64'b0000000000000000011111100000000000000000000000000000000000000000,64'b0000000000000001111000011100000000000000000000000000000000000000,64'b0000000000001111110001111100000000000000000000000000000000000000};
assign input_o[2] = {64'b0000100000000000000000000000000000000000000000000000000000000000,64'b0000100000000000000000000000000000000000000000000000000000000000,64'b0000100000000000000000000000000000000000000000000000000000000000,64'b0000100000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000001111111111,64'b0000000000000000000000000000000000000000000000000000000111111111,64'b0000000000000000000000000000000000000000000000000000000111111111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000111110000000000000000000000000000000000,64'b1111000000000000000000000001110000000000000111111111111100000000,64'b1110000000000000000000000011000000000000000000000000000000000000,64'b1111100000000000000000000011000000000000000000111000000000000000,64'b1110000000000000000000000011000000000000000001111111111110000000,64'b1100000000000000000000000001000000011000000000011100000000000000,64'b0000000000000000000000000001000000000000000110000111111100000000,64'b0000000000000000000000000000100000100000000000000111111000000000,64'b0000000000000000000000000000010000000000000000000001111100000000,64'b0000000000000000000000000000000000011000000000000001111100000000,64'b0000000000000000000000000000000000011100000000000000000000000000,64'b0000000000000000000000000000001100011100000000000000000000000000,64'b0000000000000000000000000000001100011110000000000000000000000000,64'b0000001111000000000000000000001100000010000000000000000111000000,64'b0001111111110000000000000000000011111110000000000000011111111111,64'b0000000011000000000000000000111111111111000001111111111000000001,64'b0000000011100000000000000000000000000000000111111111111000000000,64'b0000000000000000000000000000000000001111111111111111110000000000,64'b0100000000000000000001100000000011111111111110001111100000000000,64'b0000000000000000000000000000000111111111110000111111000000000000,64'b0000000000000000000011111111111111000000000000011000000000000000,64'b1111000000000000000011111111111100001111110000000000000000000000,64'b0000000000000000011110000001111111111111110000000000000000000000,64'b0000000111111111111110011111111000000000000000000000000000000000,64'b0000000001111110000000000000000000000000000000000000000000000000,64'b0000000001111110000000000000000000000000000000000000000000000000,64'b0000000011111100000000000000000000000000000000000000000000000000,64'b0000000011111000000000000000000000000000000000000000000000000000,64'b1000000010100000000000000000000000000000000000000000000000000000,64'b0000100000110000000000000000000000000000000000000000000000000000,64'b0000000000111000000000000000000000000000000000000000000000000000,64'b1000000000111000000000000000000000000000000000000000000000000000,64'b1100000000011000000000000000000000000000000000000000000000000000,64'b1100000000100000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000};
assign input_o[3] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000011111111,64'b0000000000000000000000000000000000000000000111111111111111000111,64'b0000000000000000000000000000000000000000000111111111111111111000,64'b0000000000000000000000000000000000000000000000000111111111111111,64'b0000000000000000000000000000000000000000000000000000000111111111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000011000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000010000000000000000000000000000000000,64'b0000000000000000000000000011111111111000000000000000000000000000,64'b0000000000000000000000000000000011110000000000000000000000000000,64'b0000001111111000000000000111111111110000000000000000000000000000,64'b0000000000111111110000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000100000000000000000000000000000,64'b0000001111111110010000000000000000111000000000000000000000000000,64'b0000000111111111000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000001110000000000000000000000000000,64'b0000000000000000000000000000000000110000000000000000000000000000,64'b0000000000000000000000000000110000111100000000000000000000000000,64'b0000000000000000000000000000000000001000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000001111000000000011100000000000000000,64'b0000000000000000000000000000001111111111111111111000000000000000,64'b0000000000000000000000000011111111110100000001000000000000000000,64'b0000000000000000000000000011011111110111110000000000000000000000,64'b0000000000000000000000000111010111000000000000000000000000000000,64'b0000000000000000000000000111111111011110000000000000000000000000,64'b0000000000000000000000000111111100101111000000000000000000000000,64'b0000000000001111111111101111111111111111000000000000000000000000,64'b0000000000000001111111011111111110111111100000000000000000000000,64'b0000000000000000000000011111111000111111100000000000000000000000,64'b0000000000000000000001111001111111111111100000000000000000000000,64'b0000000000000000000000011111100111111011111000000000000000000000,64'b0000000000010000000000011111000000111111110000000000000000000000,64'b0000000000000000000000110111000000011111110000000000000000000000,64'b0000000000000000001100001100000000000111100000000000000000000000,64'b0000000000000000011100011111100111011110000000000000000000000000,64'b0000000000000000000010010001100000111100000000000000000000000000,64'b0000000000000000000010010000000000000000111000000000000000000000,64'b0000000000000000011111001111000000000000001111000000000000000000,64'b0000000000000000000000000000000000000000000011111110000000000000,64'b0000000000000000000000000000000000000000000000110000000000000000,64'b0000000000000000000000000000001111111111111100000000000000000000,64'b0000000000000000000000000000001111111111111111111000000000000000,64'b0000000000000000000000000000000000000000000001110000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[4] = {64'b0000000000000000000100000000000000000000000000000000000000000000,64'b0000000000000000000011100100000000000100000000000000000000000000,64'b0000000000000000000000000000000000001110000000000000000000000000,64'b0000000000000000000000000000000000001000000000000000000000000000,64'b0000000000000000000000000000000000001000000000000000000000000000,64'b0000000000000000000000000000000111000000000000000000000000000000,64'b0000000000000000000000000000000000000000000011111100000000000000,64'b0000000000000000000000000000000000000000000011110000000000000000,64'b0000000000000000000000000000000000000110000000000000000000000000,64'b0000000000000000000000000000000000001000000000110000000000000000,64'b0000000000000000011111111111100000000000000000000000000000000000,64'b0000000000000000001101111111110000000000000000000000000000000000,64'b0000000000000000001011111111111000000000000000000000000000000000,64'b0000000000000000000001111111111000000000000000110000000000000000,64'b0000000000000000000000000011111000000000000000000000000000000000,64'b0000000000000000001111101111111100111000000000100000000000000000,64'b0000000000000000000111111111111111111001011111110000001000000000,64'b0000000000000000000011110000000000011111110000000000001100000000,64'b0000000000000000000000000000000000000011111111000000000100000000,64'b0000000000000000000000000000000000000000111111110000000000000000,64'b0000000000000000000000000000000000000000010000001100000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000110000000000000000000000000000000000000000,64'b0000000000000000000001001000000000000001110000000000000000000000,64'b0000000000000000011111111000000000000111111000000000000000000000,64'b0000000000000000001001110000000000000111110000000000000000011000,64'b0000000000000000000111110000000000000110110000000000000000000000,64'b0000000000000000000100010000000000000110110000000000000000000000,64'b0000000000000011111000000000000000000111100000000000000000000000,64'b0000000000001111111100000000000000000000100000000000000000000000,64'b0000000000011111110000000000000000000001100000000000000000000000,64'b0000000000011011000000000000000000000000000000000000000000000000,64'b1100000000011001000000000000000000000000000100000000000000000000,64'b1111100000000101111111111111111111111111110000000000000000000000,64'b1111111111111111101111111111111111111100000000000000000000000000,64'b1111111111111111111111111000000000011100000000000000000000001111,64'b1111111111111111000110111111111111111100000000000000000001111111,64'b0000000110000000001110111111111001111100000000000000000000111111,64'b0000000000000000001100000001111000011100000000000000000000000000,64'b0000000000000000000110000011011000011100000000000000000000011110,64'b0000000000000000000110000111011100011100000000000000000000000000,64'b0000000000000000000111001111011100011100000000000000000000000000,64'b0000000000000000000011001111101100001100000000000000000000000000,64'b0000000000000000000011001111011101011110000000000000000000000000,64'b0000000000000000000011000111011000100110000000000000000000001110,64'b0000000000000000000011010101011100111110000000000000000000011111,64'b0000000000000000000011010101011110111100000000000000000000111111,64'b0000000000000000000011110101011010111100000000000000000011110011,64'b0000000000000000000011110101101100111100000000000000000111000001,64'b0000000000000000000001100001101110011100000000000000000111001000,64'b0000000000000000000001100001100110001100000000000000001111000000,64'b0000000000000000000000011000110000001000000000000000001111100010,64'b0000000000000000000000011000000001111000000000000000001111101100,64'b0000000000000000000000011010000000111111100000000000000111111111,64'b0000000000000000000000011000000000000000000000000000000011100110,64'b0000000000000000000000001111111110000000000000000000000000011111,64'b0000000000000000000000000111110111000000000000000000000111111111,64'b0000000000000000000000000111111111000000000000000000001100011010,64'b0000000000000000000000000000000000000000000000000000000100011001,64'b0000000000000000000000000000000000000000000000000000001000011000,64'b0000000000000000000000000000000000000000000000000000001000011000,64'b0000000000000000000000000000000000000000000000000000011110010000,64'b0000000000000000000000000000000000000000000000000000011011010000,64'b0000000000000000000000000000000000000000000000000000011110010000};
assign input_o[5] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000011111111000000000000000000000000000000000,64'b0000000000000000000000010001111000000000000000000000000000000000,64'b0000000000000000000000000011100000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000010000000000000000000000000000000,64'b0000000000000000000000000111111100100000000000000000000000000000,64'b0000000000000000000001111110011110100000000000000000000000000000,64'b0000000000000000000001110011111001111000000000000000000000000000,64'b0000000000000000000000111110001100011000000000000000000000000000,64'b0000000000000000000000001111111000111100000000000000000000000000,64'b0000000000000000001111111110001111110000000000000000000000000000,64'b0000000000000011111100000000000111101111000000000000000000000000,64'b0000000000001111100011110000001110111111100000000000000000000000,64'b0000000000001101000000010000000111111011100000000000000000000000,64'b0000000000001100010011011000000011111010110000000000000000000000,64'b0000000000011000000000111000101111111111100000000000000000000000,64'b0000000000011000000001111000110111111111111000000000000000000000,64'b0000000000010000000001000011011111110011101000000000000000000000,64'b0000000000110000000001011011111011011111100011000000000000000000,64'b0000000000110000000000001001111111111111100011110000000000000000,64'b0000000001100000000000000000011111111000011001110000000000000000,64'b0000000001100000000000001100001111100000000000111000000000000000,64'b0000000001100000000000000100000110000000000000011111000000000000,64'b0000000001110100000000000000000000000000000000001111000000000000,64'b0000000001110100000111110001101000000000000010100011100000000000,64'b0000000001011100000000001000001000000000000000000001110000000000,64'b0000000000111100000011110000001000000000000000000000111000000000,64'b0000000000011100000011110000001000000000000000000000011000000000,64'b0000000001111100000001001010001000000000000000000000011000000000,64'b0000000001100111000000101010000000000000000000000000111000000000,64'b0000000000111011001000001010001000000000000000000001110000000000,64'b0000000000011101001000001010001000000000000000000001110000000000,64'b0000000000001100000111001010001110000000000000000111110000000000,64'b0000000000001100000001001010010100000000000001111111100000000000,64'b0000000000000100000111001010010000000000000001111110000000000000,64'b0000000000000100000000001010010000000000000001100000000000000000,64'b0000000000000100000000111010000110000000000011000000000000000000,64'b0000000000000100111110101010011100000000000011000000000000000000,64'b0000000000000011111110101011111100000000000001100000000000000000,64'b0000000000000000001111101011111110000000000001100000000000000000,64'b0000000000000000000111111111100111000000000111100000000000000000,64'b0000000000000000000000011000000110000000000110000000000000000000,64'b0000000000000000000000000000000111110000000110000000000000000000,64'b0000000000000000000000000000000111110000000110000000000000000000,64'b0000000000000000000000000000000010111100000100000000000000000000,64'b0000000000000000000000000000000000110000001100000000000000000000,64'b0000000000000000000000000000000000100000001100000000000000000000,64'b0000000000000000000000000000000000111000011100000000000000000000,64'b0000000000000000000000000000000000110000011100000000000000000000,64'b0000000000000000000000000000000000110000011100000000000000000000,64'b0000000000000000000000000000000000110000011100000000000000000000,64'b0000000000000000000000000000000000110000011100000000000000000000};
assign input_o[6] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000001110000000000000000000000,64'b0000000000000000000000000000000000000000111000000000000000000000,64'b0000000000000000000000000000000000000000011000000000000000000000,64'b0000000000000000000000000000111111110000000000000000000000000000,64'b0000000000000000000000000001111111110000011111110000000000000000,64'b0000000000000000000000000001110111111111101111111000000000000000,64'b0000000000000000000000000001111001110101101111111110000000000000,64'b0000000000000000000000000111111101111111111110001111000000000000,64'b0000000000000000000000000111100011100110111110000111000000000000,64'b0000000000000000000000000111000111000000111010000111000000000000,64'b0000000000000000000000111111110111000000111110000011000000000000,64'b0000000000000000000000111111010111000000111010011111000000000000,64'b0000000000000000000001111101111110000000111011011111000000000000,64'b0000000000000000000001111001111110000011111010111110000000000000,64'b0000000000000000000011111111111100000111100001101110000000000000,64'b0000000000000000000011100111011100001100111001111100000000000000,64'b0000000000000000000111100100111100001100110011111100000000000000,64'b0000000000000000000111111010111000000000110001110000000000000000,64'b0000000000000000001101111110111000000000110011110000000000000000,64'b0000000000000000000011111001111111111011100011110000000000000000,64'b0000000000000000000000111000000111111111111110000000000000000000,64'b0000000000000000000001111101110111110011111110000000000000000000,64'b0000000000000000000001111100000001111111111110000000000000000000,64'b0000000000000000000011110010000001100011111110000000000000000000,64'b0000000000000000000011110111001000000001111110000000000000000000,64'b0000000000000000000001100010000000000111111110000000000000000000,64'b0000000000000000000001100111001000000110011000000000000000000000,64'b0000000000000000000001110111111000000110000000000000000000000000,64'b0000000000000000000000010011011000001100000000000000000000000000,64'b0000000000000000000110110110011000011000000000000000000000000000,64'b0000000000000000000111111110011000010000000000000000000000000000,64'b0000000000000000000011111100011001110000000000000000000000000000,64'b0000000000000000000011111100111111100000000000000000000000000000,64'b0000000000000000000111011101111111000000000000000000000000000000,64'b0000000000000000000111111011110111000000000000000000000000000000,64'b0000000000000000000110110011001111000000000000000000000000000000,64'b0000000000000000000010110010001100000000000000000000000000000000,64'b0000000000000000011100100010001000000000000000000000000000000000,64'b0000000000000001111111100000010000000000000000000000000000000000,64'b0000000000000011001110000000000000000000000000000000000000000000,64'b0000000000000000111100000000000000000000000000000000000000000000,64'b0000000000000000110000000000000000000000000000000000000000000000,64'b0000000000000000000000000010000000000000000000000000000000000000,64'b0000000000000000000000000110000000000000000000000000000000000000,64'b0000000000000000000000000110000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[7] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000111000000000000000000000000000000000000000,64'b0000000000000000000000011100000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000011111000000000000000000000000000000000,64'b0000000000000000000001000011111100000000000000000000000000000000,64'b0000000000000000001110111001111000000000000000000000000000000000,64'b0000000000000000000000000111111100000000000000000000000000000000,64'b0000000000000000000011111111000000000000000000000000000000000000,64'b0000000000000000000011111100000000000000000000000000000000000000,64'b0000000000000000000010000000000000000000000000000000000000000000,64'b0000000000000000000010000000001000000000000000000000000000000000,64'b0000000000000000000000111111111111000000000000000000000000000000,64'b0000000000000000000000111111111111000000000000000000000000000000,64'b0000000000000000000010000000111111000000000000000000000000000000,64'b0000000000000000000010000001111100000000000000000000000000000000,64'b0000000000000000000010000000000000000000000000000000000000000000,64'b0000000000000000000001111110000100000000000000000000000000000000,64'b0000000000000000000000011111111100000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[8] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000110000000,64'b0000000000000000000000000000000001110000000000000000111111100000,64'b0000000000000000000000000000000011110000000000000000000000000000,64'b0000000000000000000000000000001111110000000000000000000000000000,64'b0000000000000000000000000000000000010000000000000000000000000000,64'b0000000000000000000000000000000000010000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000111110000000,64'b0000000000000000000000000000000000000000000000000000111110000000,64'b0000000000000000000000000000000000000000000000000011111001000000,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000011,64'b0000000000000000000000000000000000000000000000000000010000000111,64'b0000000000000000000000000000000000000000111000000011000000000110,64'b0000000000000000000000000000000000000000111000000000000000000011,64'b0000000000000000000000000000000000000000101000000000000000000011,64'b0000000000000000000000000000111111111000001000000000000000000001,64'b0000000000000000000000000001111111111100010000000000000000000000,64'b0000000000000000000000000011111111111111111000000000000000000000,64'b0000000000000000000000000001111111111111000000001000000000000000,64'b0000000000000000000000000011001111111110000000000000000000000000,64'b0000000000000000000000000111101001111110000000001000000000000000,64'b0000000000000000000000000111111001111110000000001000000000000000,64'b0000000000000000000000000111111001110000000000000000000000000000,64'b0000000000000000000000000111111001110000000000000000000000000000,64'b0000000000000000000000000110011001111000000000000000000000000000,64'b0000000000000000000000011111111011111000000000000000000000000000,64'b0000000000000000000000011001000010010000000000000000111111111111,64'b0000000000000000000000011001000010010000000000000000000001111111,64'b0000000000000000000000001001001000010000000000000000000001111111,64'b0000000000000000000000000001001000000000000000000000000011111110,64'b0000000000000000000000000000000000000000000000000000000011111111,64'b0000000000000000000000000000000000000000000000000000000011111110,64'b0000000000000000000000000000000000000000000000000000000011111110,64'b0000000000000000000000000000000000000000000000000000111101101111,64'b0000000000000000000000000000000000000000000000000000111111001110,64'b0000000000000000000000000000000000000000000000000001111101000111,64'b0000000000000000000000000000000000000000000000000001111100010001,64'b0000000000000000000000000000000000000000000000000001111111000001,64'b0000000000000000000000000000000000000000000000000001111111000111,64'b0000000000000000000000000000000000000000000000000001101111011100,64'b0000000000000000000000000000000000000000000000000001100111000011,64'b0000000000000000000000000000000000000000000000000001111111000010,64'b0000000000000000000000000000000000000000000000000001110111101111,64'b0000000000000000000000000000000000000000000000000111111011100001,64'b0000000000000000000000000000000000000000000000000011100111100000,64'b0000000000000000000000000000000000000000000000011111111111000000,64'b0000000000000000000000000000000000000000000000111111111111000011};
assign input_o[9] = {64'b0000000000111100000000000000000000000000011110000000000000000000,64'b0000000000011100000000000000000000011111111110000000000000000000,64'b1100000000011100000000000000000000011111111110000000000000000000,64'b1000000000011100000000000000000111111100000000000000000000000000,64'b0000000000010000000000000000000000011111100000000000000000000000,64'b0000000000010000000000000000000000000001111110000000000000000000,64'b1111111111111110000000000000000000000001111111111111000000000000,64'b1111111111111101000000000000000000000000000001111111111000000000,64'b0111111111010000000000000000000000000001111110001111111100000000,64'b1111111111010111000000000000000000000000000000111111000110000000,64'b0000001000010011000000000000000000000000000000001111110001000000,64'b0000001000011011000000000000000000000000000000000000000000000000,64'b0000000000001011000000000000000000000000000000000000000000000000,64'b0000000000001001100000000000000000000000000000000000000000000000,64'b0000000000001101000000000000000000000000000000000000000000000000,64'b0000000000001111100000000000000000000000000000000000000000000000,64'b0000000000001101000001100000010000000000000000000000000000000000,64'b0000000000010000000000011000001000000000000000000000000000000000,64'b0000000000000100010000010000000000010000000000000000000000000000,64'b0000000000000000000000011000000000000000000000000000000000000000,64'b0000000000000000100111111000111001110000000001111100000000000000,64'b0000000000000000000111011111111000000000001111111110000000000000,64'b0000000000000000000011101111111111111000001111111110000000000000,64'b0000000000000000000011111000111000111111010000001100000000000000,64'b0000000000000000000000011111111001111000000111111110000000000000,64'b0000000000000000000000000000011000000000111111100000000000000000,64'b0000000000000000000000000000011000000000000000000000000000000000,64'b0000000000000000000000000000001000000000000000111111100000000000,64'b0000000000000000000000000000000001110000001111111111110000000000,64'b0000000000000000000000000010000111110000000011111110110000000000,64'b0000000000000000000000000010011110110000000001000111010000000000,64'b0000000000000000000000001100010000001110001111111001110000000000,64'b0000000000000000000000001100001111101110001111110001111100000000,64'b0000000000000000000000001110000111011110000000111111000000000000,64'b0000000000000000000000001110000000010010111000001111110000000000,64'b0000000000000000000000001110010000001000111100000000000000000000,64'b0000000000000000000000000011000000000000000000000000000000000000,64'b0000000000000000000000000001100000000000000000000000000000000000,64'b0000000000000000000000000000110111000000000001111110000000000000,64'b0000000000000000000000000001111001000000000001111100000000000111,64'b0000000000000000000000000001111001000000000000000000000000000001,64'b0000000000000000000000000001110011111111110000000000000000000000,64'b0000000000000000000000000011110011111111110000111000000000000000,64'b0000000000000000000000000011110111000000000000000000000000000000,64'b0000000000000000000000000011110111000000000000000000000000000000,64'b0000000000000000000000000011100011000000000000000000000000000000,64'b0000000000000000000000000001100011000000000010000000000000000000,64'b0000000000000000000000000011001111111000000010000000000000000000,64'b0000000000000000000000000011001111111111110010000000000000000000,64'b0000000000000000000000000011001111011110000000000000011111100000,64'b0000000000000000000000000000111111111110000001111111111111000000,64'b0000000000000000000000000001111111111111110011111111111111110000,64'b0000000000000000000000000000100000000000000000000000010000000000,64'b0000000000000000000000000000000000000000000000000000010000000000,64'b0000000000000000000000000000000000000000000000000000000110000000,64'b0000000000000000000000000000000000000000000000000000001111110000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000001100000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000001111,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[10] = {64'b0000000000000000000000000000000000000000000000000100100000000000,64'b0000000000000000000000000000000000000000000000111000000000110000,64'b0000000000000000000000000000000000000000000000001100000000010000,64'b0000000000000000000000000000000000000000000000000111000011110001,64'b0000000000000000000000000000000000000000000000000011110111111111,64'b0000000000000000000000000000000000000000000000000001111111110000,64'b0000000000000000000000000000000000000000000000000000011111100000,64'b0000000000000000000000000000000000000000000000000000000011110000,64'b0000000000000000000000000000000000000000000000000000000000011100,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000111110000000000000000000000000000000000,64'b0000000000000000000000001111111000000000000000000000000000000100,64'b0000000000000000000000011111111000000000000000000000000000001110,64'b0000000000000000000000011111111000000000000000000000000000000111,64'b0000100000000000000000011111111000000000000000000000000000011001,64'b0000100000000000000000001111111100000000000000000000000000011111,64'b0000100000000000000000000000000000000000000000000000000000111110,64'b0000100000000000000000111111111111111000000000000000000000000001,64'b0000000000000000000111111111111111111111000000000000000000000000,64'b0011100000000000011111110011111111111111100000000000000000001000,64'b0000000000000000111100000000000111110111100000000000000000000000,64'b0000000000000001110011110000000000111011110000000000000000000000,64'b0000000000000001110000000000000000001011110000000000000000000000,64'b0000000000000001110000000000000000000011110000000000000000000000,64'b0000000000000001110000000000000000000101111000000000000000111000,64'b0000000000000000110011000000000000000111111000000000000111110000,64'b0000000000000000110111110000000000011111111000000000000110110000,64'b0000000000000000111111111000000001011011111000000000000110110000,64'b0000000000000000110101111000000001011101111000000000000110110000,64'b0000000000000000110101110000000000111101101100000000000110110000,64'b0000000000000000100101110000000001011100101100000000000111111110,64'b0000000000000000000001110000000001111100101100000000000111011111,64'b0000000000000000010000110000000000101110111100000000000011100111,64'b0000000000000000011111100000000000111110111100000000000001111100,64'b0000000000000000011100000000000000011110110110000000000000011110,64'b0000000000000000001111111000000000001111110110000000000000001110,64'b0000000000000000000011111100001111111110011111100000000000001110,64'b0000000000000000000000011110111111111110110011110000000000000110,64'b0000000000000000000000011110110110111110111111101100000000000110,64'b0000000000000000000000001111110111001110111111110000000000000011,64'b0000000000000000000000001111110011001110011110000000000000000011,64'b0000000000000000000000001110110011101110000000000000000000000010,64'b0000000000000000000000001110111011101110000000000000000000000010,64'b0000000000000000000000001110111011111110000000000000000000000010,64'b0000000000000000000000000110111011111110000000000000000000000000,64'b0000000000000000000000001111111011111100000000000000000000000000,64'b0000000000000000000000001111111011111100000000000000000000000000,64'b0000000000000000000000000111111011011100000000000000000000000000,64'b0000000000000000000000000011110010111000000000000000000000000000,64'b0000000000000000000000000011110010110000000000000000000000000000,64'b0000000000000000000000000011010100000000000000000000000000000000,64'b0000000000000000000000000000010000011110000000000000000000000000,64'b0000000000000000000000000000100001100110000000000000000000000000,64'b0000000000000000000000000000000001111110000000000000000000000000,64'b0000000000000000000000000000000000011110000000000000000000000000,64'b0000000000000000000000000000000000111111000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[11] = {64'b0000000000000000000000000000000000000000000000000000000010000000,64'b0000000000000000000000000000000000000000000000000000000011001111,64'b0000000000000000000000000000000000000000000000000000000001100011,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000100000000000001,64'b0000000000000000000000000000000000000000000000010110000000000011,64'b0000000000000000000000000000000000000000000000010000000000000100,64'b0000000000000000000000000000000000000000000000011000000010001100,64'b0000000000000000000000000000000000000000000000010000000000000000,64'b0000000000000000000000000000000000000000000000000110000000100000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000100000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000100000000000000000000000000000001111000000000000000000000000,64'b0000000110000000000000000000001111111111000000000000000000000000,64'b0000000000000000000000000000000001110010000000000000000000000000,64'b0000000000000000000000000000001111000111000000000000000000000000,64'b0000000100000000000000000000011111111111100000000000000000000000,64'b0000000000000000001111000000011111111111100000000000000000000000,64'b0000000000000000000110000001110000111001110101000100000000000000,64'b0000000000000000000110000001100000000001110000011000000000000000,64'b0000000000000000000011000001100000000001110000000000000000000000,64'b0000000000000000000000000001100000000000100000100000000000000000,64'b0000000000000000000000000001100000000000000100100000000010000000,64'b0000000000000000011100000011000000000000011100100001111111100010,64'b0000000000000000101100000110000000000010101100001111110001111110,64'b0000000000000000011100000110000000000010001110111110000000011111,64'b0000000000000000011110000110000000000010001110010000000000000111,64'b0000000000000001111111100110000000000010111010000000000000000000,64'b0000000000000000000000000010000000000010111001000000000000000000,64'b0000000000000000000011000001110000000010000000000000000000000000,64'b0000000000000000000000000000111000000110000000000000000000000000,64'b0000000000000000000000000000011111100100000000000000000000000000,64'b0000000000000000000000000000011111111110000000000000000000000000,64'b0000000000000000000000000001100111111110011111101111111100000000,64'b0000000000000000000000000001110111111100000000000000110000000000,64'b0000000000000000000000100000111111111011111111000000000000000000,64'b0000000000000000000000000000001111111111111111111111111000000010,64'b0000000000000000000000000000000000011000000000000000000000000000,64'b0000000000000000000000000000000100001100000000000000000000000000,64'b0000000000000000000000000000011110000000000000000000000000000000,64'b0000000000000000000000000000011000000000000000000000000000000000,64'b1110000000000000000000000000001111000000000000000000000000000000,64'b0110000000000000000000000000000011100000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b0001100001111000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000011100000000000000000000000000000000000000000000000,64'b0000000000000000100000000000000000000000000000000000000000000000,64'b0000000000011100000000000000000000000000000000000000000000000000,64'b0000000000000001100001110000000000000000000000000000000000000000,64'b0000000000000000000001111110000000000000000000000000000000000000,64'b0000000000000000000111011111100000000000000000000000000000000000,64'b0000000000000000000011111001111000000000000000000000000000000000};
assign input_o[12] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000111111110000000000000000000000000000000000000,64'b0000000000000000011111111111111111100000000000000000000000000000,64'b0000000000000000011111111100010100001110000000000000000000000000,64'b0000000000000000111111111111111111111000000000000000000000000000,64'b0000000000000000000010000111110001111111000000000000000000000000,64'b0000000111100000000000000000000000001111000000000000000000000000,64'b0000000011000000000000000111100000000001000000000000000000000000,64'b0000000111000000000000000000000000000000100000000000000000000000,64'b0000000000000000000000000000000000000000001000000000000000000000,64'b0000000011000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1111111000000001100000000000000000000000000000000000000000000000,64'b0000000111111111000000000000000000000000000000000000000000000000,64'b0000000000011111110000000000000000000000000000000000000000000000,64'b0000000000000000001010000000000000000000000000000000000000000000,64'b0000000000000000001100000000000000001111111100000000000000000000,64'b0000000000000000000010000000000000000111001110000000000000000000,64'b0000000000000000000000000000000000000011111100000000000000000000,64'b0000000000000000000000010000000000000000011101111000000000000000,64'b0000000000000011000000000000000000000000000000011100000001111111,64'b0000000000000000000000111111000000000000000011111110000000000000,64'b0000000000000000000000011000000000000000000000001110000000000000,64'b0000000000000000000000011100001100000000000000000000000000000000,64'b0000000000000000000000000001000000000000000000000000000000000000,64'b0000000000000000000000000000011100000000000001111100000000000011,64'b1111010000000000000000000000000000000000000011111110000000000000,64'b0011111100000000000000000000000000000000000001111001100000000000,64'b1111111100000000000000000000000000000000000000000000000000000000,64'b0000000000000111111111000000000000000000000000000000000000000000,64'b0000000000001001111111111111000000000000000000000000000000000000,64'b0000000000000011111110011111111100000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000011110000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[13] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000010000000000000000000000000,64'b0000000000000000000000000000000000000011110000000000000000000000,64'b0000000000000000000000000000000000000010100000000000000000000000,64'b0000000000000000000000000000000000000010000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000001000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000001111000000000000000000000,64'b0000000000000000000000000000000000000001111000000000000000000000,64'b0000000000000000000000000000000000000001111000000000000000000000,64'b0000000000000000000000000000000000000001101100000000000000000000,64'b0000000000000000000111111000000000000001111100000000000000000000,64'b0000000000000000011111111111111110000001111110000000000000000000,64'b0000000000000000000111111011111110011001101110000000000000000000,64'b0000000000000000011111111111111001111001011100000000000000000000,64'b0000000000000000000011111111111111111111011000000000000000000000,64'b0000000000000000000001111000000111111111111000000000000000000000,64'b0000000000000000000001110000000000111100000000000000000000000000,64'b0000000000000000000000110000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000001000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000011000000000000000000000000000000000,64'b0000000000000000000000000000110000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000100000000000000000000,64'b0000000000000000000000000000000000000000011100011110110000000000,64'b0000000000000000000000000000000000000001111100000000111100000000,64'b0000000000000000000000000000000000000111111110000000011100000000,64'b0000000000000000000000000000000001111111111110000000011110000000,64'b0000000000000000000000000000000111111110000111000000000000000000,64'b0000000000000000000000000000011111111110011111000000000000000000,64'b0000000000000000000000000000111110111111010111100000000000000000,64'b0000000000000000000000000000110001111111111111110000000000000000,64'b0000000000000000000000000000100110111111111111110000001111100000,64'b0000000000000000000000000000000000000000001101111000001100000000,64'b0000000000000000000000000000000000000010001111111000000000000000,64'b0000000000000000000000000000011111111110001111111110000000000000,64'b0000000000000000000000000000011111111110001111111000000000000000,64'b0000000000000000000000000000011110011110000011011000000000000000,64'b1111110000001110000000000000011011111100110011011000000000000000,64'b0111111101111111100000000000110000000000000111011100000000000000,64'b1111100001111110011000000000110000100000000111111100000000000000,64'b0001111110111111110000000000110000000000000111011100000000000000,64'b0001111111000011111110000000100000000000000111011100000000000000,64'b0000111011100000001111111011100001000000000111011100000000000000,64'b0000011111000000000000010000000011000000111101111100000000000000,64'b0000011111000000001111100000000111000000000111111100000000000000,64'b0000000000000001111110000011111111110000011111000000000000000000,64'b0000000011111111111100000011111111110000000000000000000000000000,64'b0000000111111111110010000000000000111000000000000000000000000000,64'b0000000111111110001111000000000000000000000000000000000000000000,64'b0011110011011111001011110000000000000000000000000000000000000011,64'b1111111111011010001011100000000000000000000000000000000000111100,64'b1111111111011010001011101100000000000000000000000000000001111100,64'b1111110110111110001011101100000000000000000000000000000001000000,64'b1101110001100010001011100000000000000000000000000000001000111000,64'b1101111011111010001011000000000000000000000000000001111000111000,64'b1111110111111001111111101111000000000000000000000000000000000000};
assign input_o[14] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000011100000000000000000,64'b0000000000000000000000000000000000000000000011100000000000000000,64'b0000000000000000000000011111100000000000000011100000000000000000,64'b0000000000000000000010000000000000000000000001000000000000000000,64'b0000000000000000000111100000000100000000000000000000000000000000,64'b0000000000000000000110100111111000000000000000010000000000000000,64'b0000000000000000010001110110111110000000000000000000000000000000,64'b0000000000000000000001111110111111100000000000000000000000000000,64'b0000000000000000000001110100101110011100000011010000000000000000,64'b0000000000000000000000010001111111110110000011010000000000000000,64'b0000000000000000111100000000111111110000000000110000000000000000,64'b0000000000000001111100000010111111000000111100000000000000000000,64'b0000000000000011111000000111100111000100110000000000000000000000,64'b0000000000000000111100000011100000000000000000000000000000000000,64'b0000000000001000000011111111110000000000000000000000000000000000,64'b0000000000001100101111100000001100111110000000000000000000000000,64'b0000000000001100100000000000000000010000000000000000000000000000,64'b0000000000001100011110000000000000000000110000000000000000000000,64'b1100000000000011100011000000000000000000110000000000000000000000,64'b0000000011100111100011100000000000000010110000000000000000000000,64'b0000000000010011100111100000000100000010110000000000000000000000,64'b0000000000100101100100000000000111000000110000000000000000000000,64'b0000000000100100111111110000000111000000011000000011111100000000,64'b0000000000111110011000000000000111000000001100000000111000001111,64'b0111111000101011110001100001111110000000000100000000000001111111,64'b0000000000111111111000000000000000000000000110000000000000000000,64'b0000000000000111111111000000000000000000000110000000000000000000,64'b0000000000000011111111111010000000000000000110000000000000000000,64'b0000000000000000001111110000000000000000000110000000000000000000,64'b0000000000000000000001111111000111111100000011000000000000000000,64'b0000000000000000000000001110000011111100001011100000000000000000,64'b0000000000000000000000001110010011110111000111100000000000000000,64'b0000000000000000000000000111000001111011110111100000000000000000,64'b0000000000000000000000000011101111111011111011110000000000000011,64'b0000000000000000000000000001100010111100111000110000000000001100,64'b0000000000000000000000000000110000111100111000110000000000000000,64'b0000000000000000000000000000111100011100011000110000000000000000,64'b0000000000000000000000000000111100011100011100111000000000000000,64'b0000000000000000000000000000011100001110001100111000000000000000,64'b0000000000000000000000000000011100001110001110111000000000000000,64'b0000000000000000000000000000000110000111000111111000000000000000,64'b0000000000000000000000000000000111000111000111111000000000000000,64'b0000000000000000000000000000000111100111000011011000000000000000,64'b0000000000000000000000000000000101100111100011011000000000000000,64'b0000000000000000000000000000000100110111100011100000000000000000,64'b0000000000000000000000000000000000111011000001110000000000000000,64'b0000000000000000000000000000000000011111000001100000000000000000,64'b0000000000000000000000000000000000001111000001001100000000000000,64'b0000000000000000000000000000000000011111000000000000000000000000,64'b0000000000000000000000000000000000000000000000011000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[15] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000011111111000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000111111111111100111100000000000000000000000001100011111,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1001100000000000000000000000000000000000000000000000000000000000,64'b1101000000000000000000000000000000000000000000000000000000000001,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000011111000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000011000000000000000000000000000000000000000000,64'b0001111111111110000001100000000000000000000000000000000000000000,64'b0011110000000000000001000000000000000000000000000000000000000000,64'b0000000000000001111111000000000000000000000000000000000000000000,64'b0000000000001111111000000000000000000000000000000000000000000000,64'b0000011111100000000000000000000000000000000000000000000000000000,64'b0000000000000001111111100000000000000000000000000000000000000000,64'b0000000111100000000011100001100101000000000000000000000000000000,64'b0000000000000000000000000000100110000000000000000000000000000000,64'b0000000000000000000000000000100111000000000000000000000000000000,64'b0000000000000000000000000011100111100000000000000000000100000000,64'b0000000000000000000000000000000111000000000000000000000100000000,64'b0000000000000000000000000000000111110000000000000000000000000000,64'b0000000000000000000000000000000110000000000000000000000000000000,64'b0000000000000000000000000000000011000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[16] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000001111111111110000000000000,64'b0000000000000000000000000011111111000011111111111111111110000000,64'b0000000000000000000000000001111110000110001000000000110111000000,64'b0000000000000000000000000011111111100011000011100000000000000000,64'b0000000000000000000000001111111110000111100000000000000000000000,64'b0000000000000000000000000011111100000011110000000000000000000000,64'b1110000000000000000000000011110000000011111111000000000000000000,64'b1101000000000000000000000000000000000000000011000000000000000000,64'b1010000000000001110000000000000000000000000001110000010000000000,64'b1111100000000011000000000000000000000000000000111001100011000000,64'b0110011111001001100100000000000000000000000000000111001100001000,64'b0000001111100111000000000000000000000000001111100111111000000000,64'b0000000001111001110000000000000000000001110000000000011111111111,64'b0000000000111110010000000000000000000000001111000000000000001001,64'b0000000000000110010000000000000000000000000000000001000000011111,64'b0000000000000111001110000000000000000000000111100001111111111110,64'b0000000000001111001111110000000000000000000000011111100000010001,64'b0000000000000011000000000000000000000000000000011111000000111001,64'b0000000000011100000000000000000000000000000001111110000000000000,64'b0000000000011000000000000000000000000000000000111100000000111001,64'b0000000000100000000000000000000000000000000000111100000000000110,64'b0000000000100100000000000000000000000000000000011111100000000110,64'b0000000000000110000000000000000000000000000000001111111111100110,64'b1111000000000110000000000000000000000000000000000000000000001000,64'b1111100000000011000000000100000000000000000000000111111100000000,64'b1111110000000010000000000100111000000000000000000000000000010000,64'b0111100000000010000000000011110000000000000000000000010000010000,64'b0000000000000110000000000000011000000000000000011111100000000000,64'b0000100000001100000000000000001100000000000000000000000001100000,64'b0000100000000111000000000000000110000000000000000000000000000000,64'b0000000000000001111000000000000011000000000000000000000000000000,64'b0000000000000000000000000000000000100000000000000000000000000000,64'b0000000000000000000000000000000000110000000000000000000000000000,64'b0000000000000000000000000000000000010000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000100000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000001000000000000000000000000,64'b0000000000000000000000000000000000000001000000000000000000000000,64'b0000000000000000000000000000000000000001000000000000000000000000,64'b0000000000000000000000000000000000000001000000000000000000000000,64'b0000000000000000000000000000000000000001000000000000000000000000,64'b0000000000000000000000000000000000000001000001010000000000000000,64'b0000000000000000000000000000000000000001000001110000000000000000,64'b0000000000000000000000000000000000000011100111110000000000000000,64'b0000000000000000000000000000000000000001011101100000000000000000,64'b0000000000000000000000000000000000000000111111100000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000001110000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[17] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000001111110000000000000000000000000000000000,64'b1100000000000000000011111111111000000000000000000000000000000000,64'b0000000000000000000011111011111110000000000000000000000000000000,64'b0000000000000000000011111111111110000000000000000000000000000000,64'b0000000000000000000011110011111111000000000000000000000000000000,64'b0000000000000000000001110111011111000000000000000000000000000000,64'b0000000000000000000000111110001111100000000000000000000000000000,64'b0000000000000000000000000111110111000000000000000000000000000000,64'b0000000000000000000000000011111111111111000000000000000000000000,64'b0000000000000000000000000001111111111111100000000000000000000000,64'b0000000000000000000000110000000000000111110000000000000000000000,64'b0000000000000000000011101110000000000111111000000000000000000000,64'b0000000000000000000000111111100000011111011000000000000000000000,64'b0000000000001111100000011101111111111111110000000000000000000000,64'b0000000010001011100000011111111111111111110000000000000000000000,64'b1111111111011110001111111100011111111110111110000000000000000000,64'b1101111111001100111111110000000000011111111000000000000000000000,64'b1100000000000111111101110000000000000000111111100000000000000000,64'b1000000000000001101111110000000000000000001111110000000000000000,64'b1000000000000000111111000000000000000000000111111000000000000000,64'b0000000000000000001111110000000000000000000001111100000000000000,64'b1000000000000000000000000000000000000000000000010111000000000000,64'b0000000000000000000000000000000000000000000000000011100000000000,64'b0000000000000000000000000000000000000000000000000001110000000000,64'b0000000000000000000001000000000000000000000000000010001111111110,64'b0000000000000000000100000000000000000000000000000010001000000111,64'b0000000000000000000110000000000000000000000000000011101111111111,64'b0000000000000000000110011001001000000000000000000000111100000001,64'b0000000000000000000101111111100100000110000000000000011000000000,64'b0000001111111111111111001111111101100111000000100000000111111111,64'b1111111100001111111111101000001110111111111111111000111111111000,64'b1111111110111111111111011000001011111100111100000000011111111111,64'b1111111110000111111111100001111111110000001111111000100101000010,64'b1011111110000000110000000000001100110000001111111100111000111000,64'b0011110000000000001000001001111111110000000110000011111110000000,64'b0000000000000000000011111111111110111000001110010001000100000000,64'b0000000000000000000001011111011111111100011011111111110101000000,64'b0000000000000000000000101111111101111100000111111111100111000111,64'b0000000000000000000111111000101111111100000000000111111101000101,64'b0000000000000000000000110111111111100000001000000001010100111111,64'b0000000000000000001111110011001000101000000000000000111101011111,64'b0000000000000011111111111111000000001000000000000000110001111100,64'b0000000000111111111111100000000101100000000000000011111111110000,64'b0000000111111111110000000000000110000000000000001111110111100000,64'b0001111101111100000000000000000000000000000000111111111110000000,64'b1111111111110000000000000000000000000000111111111101111100000000,64'b1111111000000000000000000000000000000000111111111111100000000000,64'b1111100000000000000000000000000000000000111111111110000000000000,64'b1000000000000000000000000000000000000000111111110000000000000000,64'b0000000000000000000000000000000000000000011110000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[18] = {64'b1100000000000000000000000000000000000000000000110000100000000000,64'b1100000000000000000000000000000000000000000000101000000000000000,64'b1100000000000000000000000000000000000000000000000110001110000000,64'b1100000000000000000000000000000110000000000000000111001000000000,64'b1100000000000000000000000000001100011000001100001111100000000000,64'b1100000000000000000000000000001111110000111111000001111000000000,64'b1100000000000000000000000000000001111100110111100000111000000000,64'b1100000000000000000000000000000011111111111000010000011000000000,64'b1100000000000000000000000000000000101101011000011111111110000000,64'b1100000000000000000000000000000001110001011111001101111111000000,64'b1100000000000000101000000000000000011111011001000111100011000000,64'b1100000100000000010111111111000000011111110000000000000100100000,64'b1100111100000000000000000000100000011011110001000000100001101000,64'b1111100000000001001000111100100000110011000000000000001111101000,64'b1100100001000111000000000000000000110111000000000000001100110000,64'b1100000001111101011000000000010110110111110000000000001100110000,64'b1100000001111101010000000000000000010111110000000000010111111000,64'b1100000001010001111000000000000000011110100000000000010011101000,64'b1100000000110011110000000000000001111111000000000000001000011000,64'b1100000000010111100000000000000001111011001000000000000110000000,64'b1100000000010000100000000000000001111110100000000000000000000000,64'b1100000000001100000000000000000000000000000000000000100000000000,64'b1100000000000100000000000000000000000000000000000000000000000000,64'b1100000000000100000000000000000000100000001100000000011000000000,64'b1100000000000000000000000000000000100000000000000000000000000000,64'b1100000000111110000000000000000000100000001100000000000000000000,64'b1100000000111100000000000000000000100011110000000000000011000011,64'b1100000000111000000000000000000000100010000000000000000000000000,64'b1100000000111000000000000000000000100010000000000000000000000000,64'b1100000000001100000000000000000000000010000000000000000011000000,64'b1100000001011100000000000000000000000110000000000000011000000000,64'b1100000000111110000000000000000000000110000000000000000011100000,64'b1101000000111110000000000000000000000111000000000000001001000000,64'b1100000000111100000000000000000000000011100000000000000000000000,64'b1100000000110100000000000000000000000001110110000000000000000011,64'b1100000000100110000000000000000000000000111000000000000000000000,64'b1100000000111110000000000000000000000000111000000000000000000000,64'b1100000000111110000000000000000000000000011110000000000000000000,64'b1100000000011100000000000000000000000000001110000000000000000000,64'b1100000000011100000000000000000000000000010111100000000000000000,64'b1100000000001100000000000000000000010000000011111000100000000000,64'b1100000000001111100000000000000000000100111011111111000000000000,64'b1100000000000110100000000000000000111111111001101111110000000000,64'b1100000000000111000000000000000000111111111110011111111000000000,64'b1100000000000011100000000000000000111011111000010011111000000000,64'b1100000000000001111111100100000000111101111111111111111000000100,64'b1100000000000001111110111100111111111100001111101101111000000100,64'b1100000000000001111111111111010011101110000011111110111110000100,64'b1100000000000001111111111111111100001111000001111100011110000100,64'b1100000000000000111111111011111111111011100000111111001100000100,64'b1100000000000000001111111011111111100001100000000111101100000100,64'b1100000000000000000001110000001111010101110000000001111100000100,64'b1100000000000000000000000000000011110100111000000000111100000100,64'b1100000000000000000000000000000000111111011000000000011100000000,64'b1100000000000000000000000000000000011111111100000000000000000000,64'b1100000000000000000000000000000000001111111110000000000000000000,64'b1100000000000000000000000000000000000111011111000000000000000000,64'b1100000000000000000000000000000000000111001111000000000000000000,64'b1100000000000000000000000000000000000111100011000000000000000000,64'b1100000000000000000000000000000000000011100111100000000000000000,64'b1100000000000000000000000000000000000001111111000000000000000000,64'b1100000000000000000000000000000000000000111111100000000000000000,64'b1100000000000000000000000000000000000000110000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000};
assign input_o[19] = {64'b0000000000000000011000000010100000000001100000000000000000000000,64'b0000000000000000011000000110010000000001100000000000000000000000,64'b0000000000000000001001000010001000000011100000000000000000000000,64'b0000000000000000001001000011101000000011000000000000000000000000,64'b0000000000000000000011000001101000000110000000000000000000000000,64'b0000000000000000000001100000110000111111000000000000000000000000,64'b0000000000000000000001101101111111111111100000000000000000000000,64'b0000000000000000000001110110111111100000010000000000000000000000,64'b0000000000000000000000111011111111000000000000000000000000000000,64'b0000000000000000000000011001110100000000000000000000000000000000,64'b0000000000000000000000011101111000000000000000000000000000000000,64'b0000000000000111000000000110101000000000000000000000000000000000,64'b0000000000011111100000000111101000000000000000000000000000000000,64'b0000000000111011100000000001111000000000000000000000000000000000,64'b0000000000110111100000000000000000000000000000000000000000000000,64'b0000000000110001100011100000100000000000000000000000000000000000,64'b0000000000111101110001111111100000000000000000000000000000000000,64'b0000000000111111110000000110000000000000000000000010000000000000,64'b0000000000011111100000010000000000000000000000000010000000000000,64'b0000000000001111100000000010000000000000000000000000000000000000,64'b0000000000000011000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000010000000000000000111110000000000000,64'b0000000000000000000000000000000000000000000000011110000000000000,64'b0000000000000000000000000010001000000000000000100100000000000000,64'b0000000000000000000000000010110100000000000000011101111000000000,64'b0000000000000000000000000001111010000000000000011000011000000000,64'b0000000000000000000000000000001000100000000000000001110000000000,64'b0000000000000000000000000001000010010000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000001100000000000000100000000000000000000000000000,64'b0000000000000000001111000000000000000000000000000000000000000000,64'b0000000000000000000100000000000000000000000000000000000000000000,64'b0000000000000000001100000000000000111100000000000000000000000000,64'b0000000000000000000000000000000000110000000000000000000000000000,64'b0000000000000000000000000000000011000000000000000000000000000000,64'b1100000000000000000000000000000011000000000000000000000000000000,64'b0011100000000000000000001111111111000000000000000000000000000000,64'b0000100000000000000000000000011110000000000000000000000000000000,64'b0010100000000000000000000000011000000000000000000000000000000000,64'b0000110000000000000000000111111000000000000000000000000000000000,64'b0111110000000000000000000011110000000000000000000000000000000000,64'b1110110000000000000000000001111000000000000000000000000000110000,64'b0110110000000000000000000000111100000000000000000000000000000000,64'b1111111000000000000000000000000110000000001100000000000000000000,64'b1111111000000000000000000000000110000000000110000000000000000000,64'b1111110000000000000000000000000001110000111000000000000000000000,64'b1111110000000000000000000000000000000000001000000000000000000000,64'b0000000000000000000000000000000000000000000001000000100000000000,64'b1100000000000000000000000000000000000000000000010000000000000000,64'b1110000000000000000000000000000000000000000010010001000110000000,64'b0100000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000111000000000000,64'b0000000000000000000000000000000000000000000000101111100000000000,64'b0000000000000000000000000000000000000000000000000011100000000000,64'b0000000000000000000000000000000000000000000000011111000000000000,64'b0000000000000000000000000000000000000000000000000110000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[20] = {64'b0000000000000000000000000000000000000011101000110100000111011110,64'b1111000111111000000000000000000000000011101100111100000111011110,64'b0000000111000000000000000000000000000011111110011000000111011111,64'b0000000011110000000000000000000000000011111100010100011111011111,64'b0000000011111000110000000000000000000001111110111100001111011011,64'b0000000000000000000000000000000000000001110000111100001111011000,64'b0000000000000000000000000000000000000001010000011000001111011000,64'b0000000000000000000000000000000000000001010000111100001111011000,64'b0000000000000000000000000000000000000001010001110000001111011000,64'b0000000000000000000000000000000000000001010001101100001111011000,64'b0000000000000000000000000000000000000001110001111100001111111000,64'b0000000000000000000000000000000000000001001111111110001111110000,64'b0000000000000000000000000000000000001111110001111000111111011000,64'b0000000000000000000000000001100001111111110101111111111111011000,64'b0000000000000000000000000000001111111111111110000000111111110011,64'b0000000000000000000000000000001111110111111110000011111111000000,64'b0000000000000000000001000111111110110011110110000000111111010000,64'b0000000000000000000011100000111001101111111110000011111001110000,64'b0000000000000000001111111000010011100111111100000000001111100000,64'b0000000000000000111111111000000000111110011000000111111110000000,64'b0000000000011111111000111000000000001010001001111111110000000000,64'b0000000011111111100000111100000100000011100111111001111111111100,64'b0000011111111100110101111111100000000000000000011111111110000000,64'b0001111111101111000001111001111111111111001111110000000000000000,64'b1111111100011110001111110011100011111111110111000000000000000000,64'b1111110000000000001111100011100000111111110000000000000000000000,64'b1100011100011110000001110011100000000001100000000000000000000000,64'b0011111111100011110011111101110000000000000000000000000000000000,64'b1000000000111100010011111100111000000100000000000000000000000000,64'b0000000000001110000010011100111100000010000000000000000000000000,64'b0111100000000000000010011100111000000010000000000000000000000000,64'b0000000000000000000000001100101100000110000000000000000000000000,64'b0000000011100000010000001111111000000100000000000000000000000000,64'b0000000111111100000001111111111100000110000000000000000000000000,64'b0000000010000011111100111101110000000110000000000000000000000000,64'b0000000011111111111100011111111000000110000000000000000000000000,64'b0000000011111000000000000000000000001110000000000000000000000000,64'b0000000000000000000000011000000000001110000000000000000000000000,64'b0000000000000000000000011000000001111110000000000000000000000000,64'b0000000000000000000000010000000001101110000000000000000000000000,64'b0000000000000000000000011001010001101110000000000000000000000000,64'b0000000000000000000000111010111001111110000000000000000000000000,64'b0000000000000000000000011011111001101110000000000000000000000000,64'b0000000000000000000000001111111001101110000000000000000000000000,64'b0000000000000000000000000001111001101110000000000000000000000000,64'b0000000000000000000000000001111101101110000000000000000000000000,64'b0000000000000000000000000000111011101110000000000000000000000000,64'b0000000000000000000000000000110001000011000000000000000000000000,64'b0000000000000000000000000000010000000011000000000000000000000000,64'b0000000000000000000000000000000111011110000000000000000000000000,64'b0000000000000000000000000000000001000000000000000000000000000000,64'b0000000000000000000000000000000001000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000010000000000000000000000000000,64'b0000000000000000000000000000000000111110000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[21] = {64'b0000000000000000111101111000000000000000000000000000100000000000,64'b1100000000000000111000001111000000000000000000000000100000000000,64'b0000000010000100010000011111111000100000000001100000100000000000,64'b0001111111000100000010011111111111000000000001100100100000000000,64'b0001111111000100000010110111111110000001100001100100100100000000,64'b0001111111111000000001111111110000100000010000100000100100000000,64'b0011111111111000000001111111110000000111000000011000100100000000,64'b0011111110001000000000000000000000000011100000011000100100000000,64'b1000000000001000000000000000000000000000000000000000100000000000,64'b1000000000000000000000000011111100000000000000000000000000000000,64'b0000011111111000000000000011011000000000000000000000001100000000,64'b0001111111111000000000000010010000000000000000000000000000000000,64'b0111111111110100000000000000000000000000000000000000000000000000,64'b1110000011111000000000000000000000000000000000000000111110000000,64'b1110001111111000000000000000000000000000000000000011111111100000,64'b0000001111100000000000000000000000000000000000000011111111100000,64'b0111010000000000000000000000000000000000000000000111100111000000,64'b1111111000000000000000000000000000000000000000000011111111100000,64'b0000000000000000000000000000000000100000000000000011011000010000,64'b0000000000000000000000000000000000100000000000000000100100110000,64'b0000000000000000000000000000000000110000000000000000100100011111,64'b0000000000000000000000000000000000110000000000000000011100001111,64'b0000000000000000000000000000000000110000000000000000000100000111,64'b0000000000000000000000000000000000100000000011100000000100000000,64'b0000000000000000000000000000000000100111001111111110000100000000,64'b0000000000000000000000000000000011111111111111111111110100000000,64'b0000000000000000000000000000000011001100001111111010000100000000,64'b0000000000000000000000000000000011000000001101011000000000000000,64'b0000000000000000000000000000000011000110001111111010000000000000,64'b0000000000000000000000000000000011100110001111110010000000000000,64'b0000000000000000000000000000000111111110001101111000000000000000,64'b0000000000000000000000000000000111111110001100011100000000000000,64'b0000000000000000000000000000000011111110001110011000000000000000,64'b0000000000000000000000000000000001111110001111011000000000000000,64'b0000000000000000000000000000000011001100000111111110000000000000,64'b0000000000000000000000000000011011111100000111111100000000000000,64'b0000000000000000000000000000011011011100000110111000000000000000,64'b0000000000000000000000000000000011111100000010000000000000000000,64'b0000000000000000000000000000010000111000000000000000000000000000,64'b0000000000000000000000000000000000000000000010000000000000000000,64'b0000000000000000000000000000000011100000000011111100111100000000,64'b0000000000000000000000000000000000100100000011111100111110000000,64'b0000000000000000000000000000000000100100000011101100100110000000,64'b0000000000000000000000000000000000100100000011111100100100000000,64'b0000000000000000000000000000000000000000000000011100111100000000,64'b0000000000000000000000000000000000011000000000111100011000000000,64'b0000000000000000000000000000000000001000000000011100010000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[22] = {64'b0000000000100000000000000000000000000000000000000000000000000000,64'b0000000010100000000000000000000000000000000000000000000000000000,64'b0000000000011100000000000011110000000111111111110000000000000000,64'b0000000000000000000000000000000111100011111100000000000000000000,64'b0000000000000000000000000000111111110011000000000000000000000000,64'b0000000000000000000000000000110000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000001111000000000000000000000000000000000000000,64'b0000000000000000000000011100000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000111100000000000000111000000000000000000000000000000000000000,64'b0111111111000000000100011100000000000000000000000000000000000000,64'b0100000000000000001111111110000000000000000000000000000000000000,64'b0100000000000000011111001111000000000110000000000000000000000000,64'b0000000000000000011000011111100000000000000000000000000000000000,64'b0000000000000000000000111101000110000110000000000000000000000000,64'b0000000000000000000000001111111000001100000000000000000000000000,64'b0000000000000000000000011111111111000000000000000000000000000000,64'b0000000000000000000000000000000010000000000000000000000000000000,64'b0000000000000000000010000000000000000000000000000000000000000000,64'b0000000000000000001011000000000000000000000000000000000000000000,64'b0000000000000000001011000000000000000000000000000000000000000000,64'b0000000000000000001011000000000000000000000000000000000000000000,64'b0000000000000000001011000000000000000000000000000000000000000000,64'b0000000000000000001011000000000000000000000000000000000000000000,64'b0000000000000000001011000000000000000000000000000000000000000000,64'b0000000000000000001011000000000000000000000000000000000000000000,64'b0000000000000000000011000000000000000000000000000000000000000000,64'b0000000000000000000001100000000000000000000000000000000000000000,64'b0000000000000000000101110000000000000000000000000000000000000000,64'b0000000000000000000110110000000000000000000000000000000000000000,64'b0000000000000000000011111000000000000000000000000000000000000000,64'b0000000000000000000011111000000000000000000000000000000000000000,64'b0000000000000000000011111000000000000000000000000000000000000000,64'b0000000000000000000011111100000000001111000000000000000000000000,64'b0000000000000000000111111100000001111111110000000000000000000000,64'b0000000000000000000100111010000011111111110000000000000000000000,64'b0000000000000000000001110011000011110110110000000000000000000000,64'b0000000000000000000000111101010011111110110000000000000000000000,64'b0000000000000000000010000011000110111111011000000000000000000000,64'b0000000000000000000010000001000111100000000000000000000000000011,64'b0000000000000000000000000000000000000000000111000000000000000000,64'b0000000000000000000000000000000001111001110011000000000000000010,64'b0000000000000000000000000000000010010111111111100000000000000010,64'b0000000000000000000000000000000000011100000100000000000000000000,64'b0000000000000000000000000000000000000001000011111101000000000000,64'b0000000000001111000000000000000000000101000011100011000000000000,64'b0000000000111111111111000000000000000011000011111110000000000000,64'b0000000000111000000000000000000000000000011111100000000000000000,64'b0000000000011110000000000000000000000000000111100000000000000000,64'b0000000011000000000000000000000000000011100001000000000000000000,64'b0000000000000000000000000000000000000100000000000000000000000000,64'b0000000000000000000000000000000000000100000000000000000000000000,64'b0011000000000000000000000000000000000001110000000000000000000000,64'b0010000000000000000000000000000000000001100000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000010000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[23] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000001000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000011111111000000000000000000000000000000,64'b0000000000000000000000011111111111000000000000000000000000000000,64'b0000000000000000000000001011111011000000000000000000000000000000,64'b0011111110000000000000001111111111000000000000000000000000000000,64'b0000011111000000000000000000000111000000000000000000000000000000,64'b0111111111000000000000000000000011000000000000000000000000000000,64'b0000011111110000000000000000000111010000000000000000000000000000,64'b1000000000011110000011110000000011111000000000000000000000000000,64'b0100000000000000001111111111111111111100000000000000000000000000,64'b1000000000000000001110011111111110000011111100000000000000000000,64'b1100000000000011111100000000100000000000111110000000000000000000,64'b0000000000000001111000100000000000000001011110000000000000000000,64'b0000000000000001111110000000000000000000011100000000000000000000,64'b0000000000000000001101000000000000000000111111110000000000000000,64'b0000000000000111111100000000000000000011110000000000000000000000,64'b0000000000001111111101000000000000000011100011110000000000000000,64'b0000000000001110111101000000000000000011000000010000000000000000,64'b0000000000000111110101000000000000000011000000000000000000000000,64'b0000000000000011100011000000000000000001100000000000000000000000,64'b0000000000000111110001000000000000000001100000000000000000000000,64'b0000000000000000000011000000000000000001100000000000000000000000,64'b0000000000000000000011000000000000000000100000000000000000000000,64'b0000000000000000000011000000000000000000110000000000000000000000,64'b0000000000000000000111000000000000000000111000000000000000000000,64'b1111111000000000000011000000000000000000011000000000000000000000,64'b0000000000000000000011000000000000000000010000000000000000000000,64'b0001100000000000000011000000000000000000010000000000000000000000,64'b0000000000000000000011000000000000000000010000000000000000000000,64'b0000010000000000000011000000000000000000010000000000000000000000,64'b0000110000000000000001000000001111000000010000000000000000000000,64'b0000000000000000000001100000111110000000110000000000000000000000,64'b0000000000000000000001110000100000000000110000000000000000000000,64'b0000000000000000000001110000100000000000110000000000000000000000,64'b0000000000000000000000111000000000000000000000000000000000000000,64'b0000001000000000000000011100000000000000000000000000000000000000,64'b0000000000000000000000011111001000000000000000000000000000000000,64'b0000000111100000000000000011000000000000000000000000000000000000,64'b0000000000000000000000000001000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000100000000000000000000000,64'b0000000000000000000000000000000000000000100000000000000000000000,64'b0000011000000000000000000000000000000000100000000000000000000000,64'b0000000000000000000000000000000000001111110000000000000000000000,64'b0000000000000000000000000000000000001100111000000000000000000000,64'b0000000000000000000000000000000000000111111000000000000000000000,64'b0000000000000000000000000000000000000011110000000000000000000000,64'b0000000000000000000000000000000000000001110000000000000000000000,64'b0000000000000000000000000000000000000011110000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[24] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0111100000001111100111111100000000000000000000000000000011100000,64'b0000000000000000000100000000000000000000000000000000000000000000,64'b0000000000000111110001110000000000000000000000000000000000000000,64'b0000001111111111111000111111000000000000000000000000000000100000,64'b0001111111111111111000011111111100000000000000000000000011111100,64'b1110111111111110011000011111111100000000000000000000000111111100,64'b1000100000001111111100000000000000000000000000000000000011111100,64'b1100101111111111111110000000000000000000000000000000000011111100,64'b1100001110001111110000000000000000000000000000000000000000000000,64'b1000000100000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000110010000000000000000000000,64'b0000000000000000000000000000000000000001111111111111110000000001,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000111111111111111111,64'b0000000000000000000000000000000000000000000000111111111111000000,64'b0000000000000000000000000000000000010000000000000000000000000111,64'b0000000000000000000000001111000000010000000001111111111111111111,64'b0000000000000000000000000000000000000000000001111111111111111111,64'b0000000000000000000000111111111111111000000000000000000000000000,64'b0000000000000000000000011111100000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000111111000000000000000000000000000000,64'b0000000000000000000000000000111000000000000000000000000000011111,64'b0000000000000000000000000001111111110000000000000000000000000111,64'b0000000000000000000000000000011110000000011110000000000000001111,64'b0000000000000000000000000000000000000000000000000111111111111111,64'b0000000000000000000000000000000000110000000000011111111111111110,64'b0000000000000000000000000000000011111111110011111111111111111111,64'b0000000000000000000000000000000111111111111111111011111111111111,64'b0000000000000000000000001001111111111111111111111011111111111110,64'b0000000000000000001111111111111111110001111111111000000000000000,64'b0000011111000001111111111111111110010001111111111100000000000000,64'b0000000111111111111111111111100000010000000000000000000000000000,64'b0001111111111111100110011111111111100000000000000000000000000000,64'b0011111111111110011111111111111111110000000000000000000000000000,64'b1111111000111111111100000000000000000000000000000000000000000000,64'b1111110000111111000000000000000000000000000000000000000000000000};
assign input_o[25] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000010000010000000000000000000000000000000000000000000,64'b0000000000000011000110000000000000000000000000000000000000000000,64'b0000000000000011100111000000000000000000000000000000000000000000,64'b0000000000000011100111000000000000000000000000000000000000000000,64'b0000000000000001100111000000000000000000000000000000000000000000,64'b0000000000000001111111000000000000000000000000000000000000000000,64'b0000000000000001111111000000000000000000000000000000000000000000,64'b0000000000000001111110000000000000000000000000000000000000000000,64'b0000000000000000111110000000000000000000000000000000000000000000,64'b0000000000000000011110000000000000000000000000000000000000000000,64'b0000000000000000011110000000000000000000000000000000000000000000,64'b0000000000000000111111111000000000000000000000000000000000000000,64'b0000000000000010000000000000000000000000000000000000000000000000,64'b0000000000000010000000000000000000000000000000000000000000000000,64'b0000000000000000000001000000000001110000000000000000000000000000,64'b0000000000000000000011000000000111111111111111110000000000000000,64'b0000000000000000000011001000000111111111111111111000000000000000,64'b0000000000000000001111101000000011101111111111111000000000000000,64'b0000000000000000111111000000000001111111111111100000000000000000,64'b0000000000000010011110100000000000011111111111000000000000000000,64'b0000000000000010000000100000000000000000000000000000000000000000,64'b0000000000000010000000100000000000000000000000000000000000000000,64'b0000000000000010000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000011000000000000000000000000000000,64'b0000000000000000000000000000000001100011100000000000000000000000,64'b0000000000000000000000010000000001101111111111000000000000000000,64'b0000000000000000000000000100010110110011111000000010111101111111,64'b0000000000000000000000000111111110011111110000000000000000010000,64'b0000000000000000000000000001000000000111100000000000000000000000,64'b0000000000000000000000011111111100011100000000000000000000000000,64'b0000000000000000000000011111111000011000000000000000000000000000,64'b0000000000000000000000111000000000010000000011000000000000000000,64'b0000000000000000000000111000000000110000000001100000000000000000,64'b0000000000000000000000111000000000000000000001100000000000000000,64'b0000000000000000100000011000000000000000000000111000000000000000,64'b0000000000000000000000011011000000000000011000111100000000000000,64'b0000000000000000000011110011100000000011011100000000000000000000,64'b0000000000000001111111110000000000000000001100000000000000000000,64'b0000000000000011000000000000000000000000001110000000000000000000,64'b1111111111111110000000000100000000000001101101110000000000000000,64'b0000000000000000000000000000000000000000000001111100000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000100000001110000000000000000,64'b0000000000000000000000000000000000000000000000100000010000000000,64'b0000000000000000000000000000000001111000000000000000000000000000,64'b0000000000000000000000000000000000111000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000011111,64'b0000000000000000000000000000000000000000000000000000000000011111,64'b0000000000000000000000000000000000000000000000000001111111000000,64'b0000000000000000000000000000000000000000000000001111111111011111,64'b1110000000000000000000000000000000000111111111100000011110110000,64'b1000000000000000000000000000001111111111111110000111111111110000};
assign input_o[26] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000111111000000000000000000000000000000000000000000,64'b0000000000000001111111100000000010000000000000000000000000000000,64'b0000000000000001000001100000000000000000000000000000000000000000,64'b0000000000000001000001100000000000000000000000000000000000000000,64'b0000000000000011000001000000000000000000000000000000000000000000,64'b0000000000000011000001100000000000000000000000001111111111000000,64'b0000000000000011000001100000000000000000000000001111111100000000,64'b0000000000000011000001100000000000000000000000000000000111000000,64'b0000000000000001100000000000000000000000000000000000000000000000,64'b0000000000000001100000000000000000000000000000000000000000000000,64'b0000000000000001000000000000000000000000000000000000000000000000,64'b0000000011111111000000000000000000000000000000000000000000000000,64'b1111111000011001000000000000000000000000000000000000000000000000,64'b0000001100010011000000000000000000000000000000000000000000000000,64'b0011100000000001000000000000000000000000000000000000000000000000,64'b0000000000000001000000000100000000000000000000000000000000000000,64'b0000000000000001000000000000000000000000000000000000000000000000,64'b0000000000000001000000011111000000000000000000000000000000000000,64'b0000000000000000000011110111100000000000000000000000000000000000,64'b0000000000000000000111001011100000000000000000000000000000000000,64'b0000000000000000001110001000110000000000000000000111111100000001,64'b0000000000000000001110000001110000000000000000011100001111111111,64'b0000000000000000000110001000110000000000000000111111111111111100,64'b0000000000000000000010000011100000000000000011111111110000000000,64'b0000000000000000000000000110000010000000011111100000000000000000,64'b0000000000000000000000110110001111110001111100000000000000000000,64'b0000000000000000000001111111110111111110000000000000000000000000,64'b0000000000011111000001111110111111111110000000000000000000000000,64'b0000111111111011111111111111111111110110000000000000000000000000,64'b0001111100011111111100000001110000011111111100000000000000000000,64'b0000011111111110000000010000000000011100111110000000000000000000,64'b1111111111000000000000011110110000001100011110000000000000000000,64'b1111110000000000000000011111110000000111111110000000000000000000,64'b0000000000000000000000001100110000000000111110000000000000000000,64'b0000000000000000000000001101110000000000011000111110000000000000,64'b0000000000000000000000001100110000000000011001000000000000000000,64'b0000000000000000000000000100110000000000010111111100000000000000,64'b0000000000000000000000000101110000000000000000000000000000000000,64'b0000000000000000000000000101000000000000000000000000000000000000,64'b0000000000000000000000000000000100000000000000000000000000000000,64'b0000000000000000000000000100100000000000000000000000000000000000,64'b0000000000000000000000000010011000000000000000000000000000000000,64'b0000000000000000000000000011001111110000000000000000000000000000,64'b0000000000000000000000000001100000000000000000000000000000000000,64'b0000000000000000000000000000111111111000000000000000000000000000,64'b0000000000000000000000000000011100000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000011,64'b0000000000000000000000000000000000000000000000000000000011111111,64'b0000000000000000000000000000000000000000000000000000111111111111};
assign input_o[27] = {64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100001100000000111111111100000000000000000000000000000000000000,64'b1111111111010000000000011110000000000000000000000000000000000000,64'b1100111101101000000000000100000000000000000000000000000000000000,64'b1111111111100000000000001100000001000000000000000000000000000000,64'b1111100011110000000000000000000000000000000000000000000000000000,64'b1100000001111001000000010011000000000000000000000000000000000000,64'b1110000000110110000000000001000000000000000000000000000000000000,64'b1110000000010111000000000001001000000000000000000000000000000000,64'b1101000000000001100000000000101000000000000000000000000000000000,64'b1100000000011110100011111100100000000000000000000000000000000000,64'b1100000110011110000000000000110000000000000000000000000000000000,64'b1100000111110011100000000000110000000000000000000000000000000000,64'b1100001111110011110000000000010000000000000000000000000000000000,64'b1100001100000000000000000000001100000000000000000000000000000000,64'b1100000010011100000000000000000011000000000000000000000000000000,64'b1100000000011000110000000000000011000000000000000000000000000000,64'b1100000000001000000000000000000001100000000000000000000000000000,64'b1100000000000000000000000000000000110000000000000000000000000000,64'b1100000000000000000000000000000000011000000000000000000000000000,64'b1100001100000000000000000000000000001000000000000000000000000000,64'b1100011100100000000000000000000000000100000000000000000000000000,64'b1100001111110000000000000000000000000000000000000000000000000000,64'b1110001101010000000000000000000000000001100000000000000000000000,64'b1100000101100000000000000000000000000000110000000000000000000000,64'b1100000011110100000000000000000000000000000000000000000000000000,64'b1100000000111010000010100000000010000000000110000000000000000000,64'b1100000000011001100011011111000000000000000000100000000000000000,64'b1100000000001110011111111111011000000000001110001110000000000000,64'b1100000000000111111111100011110000000000011110111110110000000000,64'b1100000000000011111111001101111000000000001101110111100000000000,64'b1110000000000000001111000000001111100000000111111001110000000000,64'b1110000000000000000000000000000000111110000001110000110000000000,64'b1111100000000000000000000000000000111110110001111011110000000000,64'b1111111000000000000000000000000000111111100000111111111000000000,64'b1100111100000000000000000000000000101111100000000001111000000000,64'b1110001100000000000000000000000000101111100000011100010000000000,64'b1100001110000000000000000000000000001001100110000000110000000000,64'b1100000110000000000000000000000000001101100000000000000000000000,64'b1100000011100000000000000000000000001101100000000000000000000000,64'b1100000001100000000000000000000000001101100000000000000000000000,64'b1100000000110000000000000000000000000111100000000000000000000000,64'b1100000000110000000000000000000000000011100000000000000000000000,64'b1100000000011000000000000000000000000000000000000000000000000000,64'b1100000000010000000000000000000000000011110000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000001110000000000000000000000000000000000000,64'b1110000000000000000000001111000000000000000000000000000000000000};
assign input_o[28] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000111000000000000000000000000000000000000000000000,64'b0000000000000000000000011110000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000001111111111000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000001111110000000000000000000000000000000000000,64'b0000000000000000000111111111000000000000000000000000000000000000,64'b0000000000000000000000110111111100000000000000000000000000000000,64'b0000000000000000000001111111000000000000000000000000000000000000,64'b0000000000000000000000111111110000000000000000000000000000000000,64'b0000000000000000000000011111110000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000001000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000111000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000111000000000000000000000000000000000000000000000000,64'b0000000000010000000000000000000000010000000000000000000000000000,64'b0000000110000000000000000000000001100000000000000000000000000000,64'b0001111000000000000000000000000001111000000000000000000000000000,64'b0000000000000000000000000000000111111000000000000000000000000000,64'b1100000000000000000000000000000111110000000000000000000000000000,64'b0000000000000000000000000000000001111111111110000000000000000000,64'b0000000000000000000000000000000000011111110000000000000000000000,64'b0000000000000000000000000000011111110001111110000000000000000000,64'b0000000000000000000000000000001111111110000000000000000000000000,64'b0000000000000000000000000000000000001111111111000000000000000000,64'b0000000000000000000000000000000111111101111111000000000000000000,64'b0000000000000000000000000000000011111111000001000000000000000000,64'b0000000000000000000000000000000000000000011110000000000000000000,64'b0000000000000000000000000000001111111000000000000000000000000000,64'b0000000000000000000000000000111111110000000000000000000000000000,64'b0000000000000000000000000000000001110000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[29] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000100000000000000000000000000000000000000,64'b0000000000000000000000001111100000000000000000000000000000000000,64'b0000000000000000000000111111111110000000000000000000000000000000,64'b0000000000000000000111111101111111111110000000000000000000000000,64'b0000000000000000111111001001111111111110000000000000000000000000,64'b0000000000000111111101111111101111100111000000000000000000000000,64'b0000000000001111111111111111111111001111100000000000000000000000,64'b0000000000011101111100011111111111100110110000000000000000000000,64'b0000000000010111110000001111111111110101111100000000000000000000,64'b0000000000010001000000000111110101111110101110000000000000000000,64'b0000000000110000000000000001110111111100001110000000000000000000,64'b0000000000110000000000000000101111111110011110000000000000000000,64'b0000000000110000010000000000011111111111001110000000000000000000,64'b0000000000110000111100000000011111111111111110000000000000000000,64'b0000000000110000001110000000000000111111111100000000000000000000,64'b0000000000110000000111110000000000011111111000000000000000000000,64'b0000000000110001011011110000000000001111111110000000000000000000,64'b0000000000110001011100111000000100000111111110000000000000000000,64'b0000000000011101001110111000000000000011111111000000000000000000,64'b0000000000001101000111100000000000000011111111100000000000000000,64'b0000000000001100010011110000000000000001111111000000000000000000,64'b0000000000001100110001100000000000001110001111000000000000000000,64'b0000000000001101011000000000000000000110001111000000000000000000,64'b0000000000001110011100000000000000000100000000000000000000000000,64'b0000000000000110001100000000000000000000000000000000000000000000,64'b0000000000000110001110000000000000000000000000000000000000000000,64'b0000000000000000001011000000000000000000000000000000000000000000,64'b0000000000000001000011000000000000001000111000000000000000000000,64'b0000000000000001000011100000000000001000000000000000000000000000,64'b0000000000000001000001110000000000000000000000000000000000000000,64'b0000000000000001000001110001111100000000000000000000000000000000,64'b0000000000000011000000110111110000001100000000000000000000000000,64'b0000000000000011000001111111110000111100000000000000000000000000,64'b0000000000000011000001111111110001111110000000000000000000000000,64'b0000000000000011000000110111011111110011000000000000000000000000,64'b0000000000000100000000000110011111111111000000000000000000000000,64'b0000000000000100000000000000010000110011000000000000000000000000,64'b0000000000001100000000000000010011100111000000000000000000000000,64'b0000000000001110000000000000000010000011110000000000000000000000,64'b0000000000001110000000000000000010000001111000000000000000000000,64'b0000000000000110000000000000000000000000001100000000000000000000,64'b0000000000000110000011110000000000000000000100000000000000000000,64'b0000000000000111000111110000000011000000000100000000000000000000,64'b0000000000000011000110110111111111000000000011100000000000000000,64'b0000000000000011111111100011111111000000000001110000000000000000,64'b0000000000000011111111000001111111000000000000011000000000000000,64'b0000000000000001111111000000001111111000000000011110010000000000,64'b0000000000000001111111000000000001111111000000000111010000000000,64'b0000000000000000111110000000000001100111010000000111000000000000,64'b0000000000000000011100000000000000000011110000000011100000000000,64'b0000000000000000000000000000000000000001110000000001100000000000};
assign input_o[30] = {64'b0110000110000000000000000000000000000000000000000000000000000000,64'b1110000100000000000000000000000000000000000000000000000000000000,64'b1100001100000000000000000000000000000000000000000000000000000000,64'b1001110000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0011000000000000000000000000000000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000001100000000000000000000000000000000000,64'b0000000000000000000000000011110000000000000000000000000000000000,64'b0000000000000000000000100111111000000000000000000000000000000000,64'b0000000000000000001100111111111100000000000000000000000000000000,64'b0000000000000000000111101100000110000000000000000000000000000000,64'b0000000000000000000100001110000110000000000000000000000000000000,64'b0000000000000000000101101111000110000000000000000000000000000000,64'b0000000000000001111111111111000111000000000000000000000000000000,64'b0000000000000001100011111101000011000000000000000000000000000000,64'b0000000000000001100001111100000011000000000000000000000000000000,64'b0000000000000001100000000000000011000000000000000000000000000000,64'b0000000000000001000000000000000001101100000000000000000000000000,64'b0000000000000011111111000000000001110010000000000000000000000000,64'b0000000000000000111111000000000000111000000000000000000000000000,64'b0000000000000000011111100000000000111100000000000000000000000000,64'b0000000000000000011011111110000000011011100000000000000000000000,64'b0000000000000000011001111100000000010011000000000000000000000000,64'b0000000000000000001110011100001000000011100000000000000000000000,64'b0000000000000000000111011100000000111111110000000000000000000000,64'b0000000000000000000011101001000000111010000000000000000000000000,64'b0000000000000000000000100100001111111111100000000000000000000000,64'b0000000000000000000000000001110001111000000000000000000000000000,64'b0000000000000000000000000000111111111000000000000000000000000000,64'b0000000000000000000000001111111111001100000000000000000000000000,64'b0000000000000000000000000111111111110000000000000000000000000000,64'b0000000000000000000000000000110111111000000000000000000000000000,64'b0000000000000000000000000001101001110000000000000000000000000000,64'b0000000000000000000000000000111010000000000000000000000000000000,64'b0000000000000000000000000001111110000000000000000000000000000000,64'b0000000000000000000000000000011110000000000000000000000000000000,64'b0000000000000000000000000000110110000000000000000000000000000000,64'b0000000000000000000000000000110110000000000000000000000000000000,64'b0000000000000000000000000000111110000000000111000000000000000000,64'b0000000000000000000000000000011100000000000001100000000000000000,64'b0000000000000000000000000000011100100000000011100000000000000000,64'b0000000000000000000000000000000000000000000010110000000000000000,64'b0000000000000000000000000000000001000000000000011000000000000000,64'b0000000000000000000000000000000000000000000010011000000000000000,64'b0000000000000000000000000000000000000000000010000000000000000000,64'b0000000000000000000000000000000000000000000001110000000000000000,64'b0000000000000000000000000000000000000000000000110000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000};
assign input_o[31] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000111100000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000011111100000000000000000000000000,64'b0000000000000000000000000000001111111100000000000000000000000000,64'b0111111000000000000000000000001111110000000000000000000000000000,64'b1111111111000000000001111100011111111000000000000000000000000000,64'b1100111111100011100001110100011111100000000000000000000000000000,64'b1111111111111100000111111100000000000000000000000000000000000000,64'b0011111111111110000111111100000000000000000000000000000000000000,64'b0011111111101100000011111100000110000000000000000000000000000000,64'b0111111111111111000000000000000000000000000000000000000000000000,64'b0001111111111110000000000000000000000000000000000000000000000000,64'b0000000111100000000011111100000000000000000000000000000000000000,64'b0000000000000111111111111111111000000000000000000001111111111111,64'b0000011111111111111111111111110000000000000000000000000111111110,64'b0011111111111111111111111111110000000000000000000001111111111111,64'b0001111111111011111111111100110000000000000000000011111111111111,64'b0000111111001111111111111000000000000100000000000000000111111111,64'b1111100111111111111100111110000000000100000000000000000000000000,64'b1111011111111110000000010010000000000100000000000000000001111001,64'b1111111111111000000000000000000000000100000000000001111111111111,64'b1111111000000001111110000000000000000100000000000000000000000011,64'b1111100000000011111010000000000000000100000000000000000000000010,64'b0000000001111101110010000000000000000100000000000000000001000010,64'b1111111111111000000000000000000000000100000000000000000000000000,64'b1111111110000000000000000001100000000000000000000001111000000001,64'b1111111000001000000000000001100000000000000000000000000000000000,64'b0111110000001000000000000001100000000000000000000000000000000000,64'b1111111110000000000000000010010000000000000000000000000000001110,64'b0000000000000000000000000000000000000000000000000000000001111111,64'b0000000000000000000100000000000000000000000000000000000111111111,64'b0000000000000000100000000000000000000000000000000000000000001101};
assign input_o[32] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000011111111000000000000000000000000000000,64'b0000000000000000000000000010111111000000000000000000000000000000,64'b0000000000000000000000000011111000000000000000000000000000000000,64'b0000000000000000000000000000000000011100000000000000000000000000,64'b0000000000000000000000000000000000001110000000000000000000000000,64'b0000000000000000000000000000000000000100000011111000000000000000,64'b0000000000000000000000000010111000000011100000000000000000000000,64'b0000000000000000000000000011111100000011100000000000000000000000,64'b0000000000000000000000000011000000000000001000000000000000000000,64'b0000000000000000000000000011000000000000011100000000000000000000,64'b0000000000000000000000001101110000000111000000100000000000000000,64'b0000000000000000000000000010111111100000011111110000000000000000,64'b0000000000000000000000000010111000000000000001110000101100001110,64'b0000000000000000000000000000111000000000000000110000000000000000,64'b0000000000000000000000000000110000000000001111111111111111111111,64'b0000000000000000000000000001110000000000000111110000000001111111,64'b0000000000000000000000000001111111000100011111000000000000000000,64'b0000001111000000000000000001110010111100110000000000000000000000,64'b0000000000000000000000000000111110111101110000000000000011110000,64'b0000011111111000000000000000110011111001100000000000000000000000,64'b0001111111110000000000000001110001011110000000000000000000000000,64'b0000000000000000000000000001110011111111000000000000000000000000,64'b0000000000000000000000000000110001110111100000000000000000000000,64'b0000000000000000000000000111100111111111000000000000000000000000,64'b0000000000000000000000001111110111111111100000000000000000000000,64'b0000000000000000000000001111111111111111100000000000000000000000,64'b0000000000000000000000000111111110101111100000000000000000000000,64'b0000000000000000000000000111110001001111110000000000000000000000,64'b0000000000000000000000000001111001101110100000000000000000000000,64'b0000000000000000000000000000010010111101000000000000000000000000,64'b0000000000000000000000000000110010111000000000000000000000000000,64'b0000000000000000000000000000001111011100000000000000000000000000,64'b0000000000000000000000000000000111101000000000000000000000000000,64'b0000000000000000000000000000000011110000011000000000000000000000,64'b0000000000000000000000000000000000111100011100000000000000000000,64'b0000000000000000000000000000000000111101111111110000000000000000,64'b0000000000000000000000000000000001110111111111100000000000000000,64'b0000000000000000000000000000000000101011110000000000000000000000,64'b0000000000000000000000000000000001111111110000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[33] = {64'b0000000000000000000000000010000000000000000010000000000000000000,64'b1110000000000000000000000110000000000000001011111111111111111111,64'b0011111111000000000001100110000000000000000000000000000000000111,64'b0000000000000000000000000000001000000000001000000000000000000001,64'b0000000000000000000000000001111100000000001110011111100001111111,64'b1111100000000000000111100000100000000000000000000000000001111110,64'b1111111111111111111111111111111100000000000000000000000000111111,64'b1111111111111111111111111111111100000001111111111111111111111111,64'b0000000000000000000000000000111000000111111111111111111111111111,64'b0000000000000000000000000000000000111111111111111111111111000000,64'b0000000000000000000000000000000000011000000000111000000000000000,64'b0000000000000000000000000000000001011100001111111111100000000000,64'b0000000000000000000000011111111110000111110000000011111000000000,64'b0011111100000000000000111111111110000000000000000000000000000000,64'b0000000000000000000000111111111110000000001111111111111100000000,64'b0000000000000000000000001111111001000000000000000000000000000000,64'b0000100000000000000000001111100000000000001111111111111110000000,64'b0000000000000000000000001111000111111000000000000000000000000000,64'b0000000000000000000000000011111110000100000000000000000000000000,64'b0000000000000000000000000000111100000100000000000000000000000000,64'b0000000000000000000000000000000000000100000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000110000001111110000000000000000000000000,64'b0000000000000000000000000000000011100000000000000000000000000000,64'b0000000000000000000000000000000000110000000000000000000000000000,64'b0000000000000000000000000000000000100000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000001110000000000000000000,64'b0000000000000000000000000000000000000000001111000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000001011100000000000000000000000000000000000000,64'b0000000000000000000000001111000000000000000000000000000000000000,64'b0000000000000000000000011100000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000011100000000000000000000000000000,64'b0000000000000000000000000000000000100000000000000000000000000000,64'b0000000000000000000000000000011100110000000000000000000000000000,64'b0000000000000000000000000000000011100000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000011100000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000111000010000000000000000000000000,64'b0000000000000000000000000000001111111000000000000000000000000000,64'b0000000000000000000000000000000111111111110000000000000000000000,64'b0000000000000000000000000000000111111000000000000000000000000000,64'b0000000000000000000000000000000000111111100000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000111111111111111000000000000};
assign input_o[34] = {64'b1111000000000000000000000000000000000000000000000010001000000000,64'b1110000111111000001000100000000000000000000000000010001000000000,64'b1111000000001000001000000000000000000110010000000010001000000000,64'b1100000000000000000000000000000000000110010000000000001000000000,64'b0000000000000000000000000000000000000110010000000000001000000000,64'b0000000000000000000000000000000000000110010000000000001000000000,64'b0000000000000000000000000000000000000110010000000000111000000000,64'b0000000000000000001000000000000000000010010000000001111000000000,64'b0000000000000000001000000000000000000011010000000001111000000000,64'b0000000000000000001000000000000000000010010000000001111000000000,64'b0000000000000000001000000000000000000010010000000001111000000000,64'b0000000000000000111100000000000000000010000000000001110010000000,64'b0000000000000001111111000000000000000001000000000000011010000000,64'b0000000000000001110110000000000000000000000000000000001100000001,64'b0000000000000000110111000000000000000000000000000000000100000001,64'b0000000000000000001011000000000000000000000000000000000000000000,64'b0000000000000000001011000000000000000001110000000000000000000000,64'b0000000000000000001011000000000000000000000000000000000000000000,64'b0000000111111000001011000000000000000000010000000000000000000000,64'b0000000111110000111111000000000000000000100000000000000000000000,64'b0000000011100001110111000000000000000001111000001100000000000000,64'b0000000000000001111011000000000111000001111111111111100000000000,64'b0000000000000001110011000000000000000000000011100011100000000000,64'b0000000000000001111111000000000000000000000011110111000000000000,64'b0000000000000011001001000000000000000000000011110111000000000000,64'b0000000000000000011100110000000000000000000001110111000000000000,64'b0000000000000001111100110000000000000000000000110011000000000000,64'b0000000000000011111010110000000000000000000000011011000000000000,64'b0000000000001110000110111000000000000000000000011001000000000000,64'b0000000000001000000110111000000000000000000000010001000000000000,64'b0000000000000001111111111000000000000000000011111100011111111000,64'b0000000000000011111111110000000000000000000001111100111111111000,64'b0000000000000011001101110000000000000011110111110111111111000001,64'b0000000000000000001101110000000000011001111111111111111101111111,64'b0000000001110000001011110111100011111000000000111111111111111110,64'b0000000111111001000111101111111111111100000000111111111111100000,64'b0000000001001111111111111111111011111100000000011111111111000000,64'b0000001111111111111111111111111111111100000000000011100000000000,64'b0000001011110000001111111111111011111000000000000000000000000000,64'b0000111111111111100000001111111111101100000000000000000000000000,64'b0000011000111111100000001111111111111110000000000000000000000000,64'b0000001000000000000000011111110001111110000000000000000000000000,64'b1111111000000000000000001110110000111011000000000000000000000000,64'b0111111111111111111111111100110000111011000000000000000000000000,64'b0000011111111111111111111000010001111001000000000000000000000000,64'b0000001111111111111111111000010001100110000000000000000000000000,64'b0000001111110111111111100000000000001111100000000000000000000000,64'b0000001011111111111111100000000000111111111100000000000000000000,64'b1111111101111111111111100000000001111111111000000000000000000000,64'b1111111111111111111111111111111100000000000000000000000000000000,64'b1111111111111100000000000000000000000000000000000000000000000000,64'b1111111111110000000000000011111111111111100000000000000000000000,64'b1111111100000000000000000000000000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000011110000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[35] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000011,64'b0000000000000000000000000000000000000000000011111111000000000010,64'b0000000000000000000000000000000000000000000011111111100000000011,64'b0000000000000000000000000000000000000000000001111001100000011111,64'b0000000000000000000000001000000100000000010000000000110001111111,64'b0000000000000000000000001000100100000000011000000000111000001111,64'b0000000000000000000000001000100100000000111100000000111000000001,64'b0000000000001000000000001000000000000000011101000011111100000000,64'b0000000011111111111111111100011000000000011100000010111100000000,64'b0000000000001000000001111111111111111110011111000011111100000000,64'b0000000000001111111111111011111100000000011110000011111000000000,64'b0000000011111111111111111111111100000000001111000011111000000000,64'b0000000011111111111000000111111100000000000111100010111000000000,64'b1111111111111111111110000011111100000000000011100010111000000000,64'b1111110000000000011110000011111100000000000011100110111000000000,64'b0000000000000000011110000011111100000000000011100100111000000000,64'b0000000000000000011110000011111000000000000011100100111000000000,64'b0000000000000000001110000011111100000000000001111011111000000000,64'b0000001110000011101110001011011100000000000000011110110000000000,64'b1111111111111000001110001111011100000000000000011111000000000000,64'b1111111000000000001110001111011100000000000000000111000000000000,64'b0000000000000000001110001000011000000000000000000010000000000000,64'b0000000000000000001110000000010000000000000000000000000000000000,64'b0000000000000000001110000000000011100000000000000000000001111111,64'b0000000000000000000110000000000011110000000000000000000001111111,64'b0000000000000000000000010100000000000000000000000000000000111111,64'b0000000000000000000000111100000011111100000000000000000000111111,64'b0000000000000000000000011111111111111100000000000000000011111111,64'b0000000000000000000000000000000000000001111000000000000000000000,64'b0000000000000000000000000000000011111111111100000000000000000000,64'b0000000000000000000000000000000011111111111000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000001111111111000000000000000000000,64'b0000000000000000000000000000000000111111000000000000000111110000,64'b0000000000000000000000000000000000000000000000000000111111110000,64'b0000000000000000000000000000000000000000000000000000111111100011,64'b0000000000000000000000000000000000000100000000000000111111111111,64'b0000000000000000000000000000000000000000000000000000011111111110,64'b0000000000000000000000000000000000000000000000000000011111110000,64'b0000000000000000000000000000000000001111000001111100100000000000,64'b0000000000000000000000001000000000001100011110000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000001111000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000011111111111111111100000000000000000000000000};
assign input_o[36] = {64'b0000000000000000000000000000000000000000000000000000011001111100,64'b0000000000000000000000000000000000000000000000000000011001111100,64'b0000000000000000000000000000000000000000000000000000011001111100,64'b0000000000000000000000000000000000000000000000000000011001111100,64'b0000000000000000000000000000000000000000000000000000011001111110,64'b0000000000000000000000000000000000000000000000000000011001111100,64'b0000000000000000000000000000000000000000000000000000011001111100,64'b0000000000000000000000000000000000000000000000000000011000111100,64'b0000000000000000000000000000000000000000000000000000011001111111,64'b1100000000000000000000000000000000000000000000000000011101111011,64'b1111100000000000000000000000000000000000000000000000011111111000,64'b1111111000000000000000000000000000000000000000000000111101111111,64'b1111111100000000000000000011110000000000000000000000111001111111,64'b1110111111111000000000111111111100000000000000000000011111111111,64'b1111111000000000000011111111111110000000000000000000011110111011,64'b1111110000010000001111111111111110000000000000000000111011111111,64'b1111111000010000001111111111011111111000000000000000111101111111,64'b0011110000011000001111111111111111111111000000000000111001111110,64'b0000000001111100001110001111111111101111000000000000011101110110,64'b0000000111111110001110000000110011111111100000000000111001111110,64'b0000000011011110000111111000111111111111100000000000111101111111,64'b0000000111111111000001101111111111111111100000000000111101111101,64'b0000000011110111000000000011111111111100110000000000111001111111,64'b0000000000111111000000001111111110000001111000000000111001111110,64'b0000000000011011100000000011111110000010111000000000111001111011,64'b0000000000011011110000000000000110000000111000000000111001111110,64'b0000000000011111111000000000111111100000111000000000111000111110,64'b0000000000001111111000000011111111111110111100000000111000111110,64'b0000000000000011111100000011111001000000011110000000111000111100,64'b0000000000000001111100000011111111100000001110000000111000111100,64'b1100000000000001001110000011111000000000000110000000111000111011,64'b1000000000000000011111000010011010000000110110000000011000111000,64'b1111100001111111111111000000011000000000110110000000011000111000,64'b1011111111111111101111100000011001000000100110000000111000111100,64'b1111111000110111111111100000011111100000001110000000011000111111,64'b0110000011111111111011111000011111100000001110000000011001111001,64'b1111100000000100000011111110010111000000001110000000011000111000,64'b0000000000000000000000011110010111000000111110000000111000111000,64'b0000000000000001000000111100001111000000111111100000111000111000,64'b0000000000000000000000111111000111000001111111100000111011011100,64'b0000000000000000000000111111000111010000011111000000111001011100,64'b0000000000000000000001111111100111001111111110000000111000111100,64'b0000000000000000000001111011110111110111111000000000111001101100,64'b0000000000110000000000000000110011111111000000000000111110011000,64'b0000000011110000000000000000010011111111000000000000111111110111,64'b1111111100010000000000011000010001110111000000000000111111111111,64'b1111111111111100000011100000010001110110000000000000111011101111,64'b0000000111110000000000000010000000110110000000000000111111101111,64'b0000000000000000000000000000000000110100000000000000111111100111,64'b0000000001111111111111100000000000110100000000000000111111101111,64'b1000111111111111111111111111111000110100000000000000111101111111,64'b1111111111111111111111111111111100110100000000000000111101100111,64'b1111111111110001111111111111111111001100000000000000111111101111,64'b0111111111111000001000011000011110000000000000000000111111100110,64'b0000000000000000000000000001011110000000000000000000111111101110,64'b0000000000000000000000000001101110000000000000000000111011101111,64'b0000000000000000000000000000111111000000000000000000111011100111,64'b0000000000000000000000000001111111000000000000000000111011100111,64'b0000000000000000000000000000011111000000000000000000111011100110,64'b0000000000000000000000000000011111000000000000000000111011100110,64'b0000000000000000000000000000011111000000000000000000111011101110,64'b0000000000000000000000000000011111000000000000000000111011100110,64'b0000000000000000000000000000011111000000000000000000111011100110,64'b0000000000000000000000000000011111000000000000000000111011100110};
assign input_o[37] = {64'b0000000000000000000000000000000000100000000000000000000000000000,64'b0000000000000000000000000000000000001111111111111111110000000000,64'b0000000000000000000000000000000000001111111111111111110000000000,64'b0000000000000000000000000000000000000000000000000000000000000100,64'b0000000000000000000000000000000000000000000000000111100000000000,64'b0000000000000000000000000000000000000000000000011111111100000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000111111000001100,64'b0000000000000000000000000000000000000000000000011111111100001111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000100000000000000000000000000000000,64'b0000000000000000000000000000000100000000000000000000000000000000,64'b0000000000000000000000000000000111110000000000000000000000000000,64'b0000000000000000000000000000000111111110000000000000000000000000,64'b0000000000000000000000000000000000111100000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000001000000000000000000000000000000000000,64'b0000000000000000000000001111000000000000000000000000000000000000,64'b0000000000000000000000000010000000000000000000000000000000000000,64'b0000000000000000000000011111000000000000000000000000000000000000,64'b0000000000000000000000011110000010000000000000000000000000000000,64'b0000000000000000000000000000000111000000000000000000000000000000,64'b0000000000000000000000000000000111000000000000000000000000000000,64'b0000000000000000000011111100001011000000000000000000000000000000,64'b0000000000000000000000011111111000000000000000000000000000000000,64'b0000000000000000000000000011100000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000001100000000000000000000000000000000,64'b0000000000000000000000001111000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000100000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000111111111110000000000001111100000000,64'b0000000000000000000000000011111111111111111111111111111111111111,64'b0000000000011111000000000000000011111111111111111000111111111111,64'b0000000000000011111100000000000000000000000000000000000000000000,64'b0000000000000011111100000000000000000000000000000000000000000000,64'b0000000000000000111110000000000000000000000000000000000000000000,64'b0000000000000000000111110000000000000000000000000000000000000000,64'b0000000000000111100011111000000000000000000000000011111111111000,64'b0000000000000000000000000000011111000000000000000000000000000000,64'b0000000000000000000000000000111111100000000000000000000000000000,64'b0000000000000000000011100001111000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000001111100000000000000000000000000000000,64'b0000000000000000000000000001111000000000000000000000000000000000,64'b0000000000000000000000000000000000000011111100000000000000000000};
assign input_o[38] = {64'b0000000000000000000000000000000000000000001100000000000000000110,64'b0000000000000000000000000000000000000000001100000000100000001110,64'b0000000000000000000000000000000000000000000110000000001111110111,64'b0000000000000000000000000000000000000000000110000001000001100111,64'b0000000000000000000000000000000000000000000110000000000000101111,64'b0000000000000000000000000000000000000000000101000000000000001110,64'b0000000000000000000000000000000000000000000011100000000000001110,64'b0000000000000000000000000000000001111111111001101000000000000111,64'b0000000000000000000000001111111000000001111111101100000000001111,64'b0000000000000000000000001111111111111111111111011110000000000011,64'b0000000000000000000000010001110000000110000111011111100000001111,64'b1000000000000000000000000111111100000111111000000011111100000000,64'b0000000000000000000111111110011000000000000011111001000000000011,64'b0000011100000000000011111111110000000000000011111111111111011111,64'b1000000000000000000001111111111111110000001111000000010111111000,64'b0000011100000000001111111111111111111111101111111111111110000000,64'b0000000000000000000000000111111111111010111111111111111100000000,64'b0000000000000000000000000000111100111000100000111100001000000000,64'b0000000000000000000000000000100111110000001111111100000000000000,64'b0000000000000000000000000000001011111000000011000000000000000000,64'b0000000000000000000000000000000000000111111111111000000000000001,64'b0000000000000000000000000010000011110000000111111100000000000111,64'b0000000000000000000000000000000111111111111111111111111000111111,64'b0000000000000000000000000100000100000000011000011111011111111110,64'b0000000000000000000000000100000100000000001100011011111111111100,64'b0000000000000000000000000100000100000000000000111000000111111100,64'b0000000000000000000000000000000111110000111101010000000010011111,64'b0000000000000000000000000000000110000000011111000000000000001111,64'b0000000000000000000000000000000111111001111111110000000000000001,64'b0000000000000000000000000000000000000111111100000000000000010000,64'b0000000000000000000000000000011111000000000100000000000000001111,64'b0000001000000000000000000011100011000111000001000000000000010000,64'b0000000000000000000000000011101011111110000000000000000000000111,64'b0000000000000000000010000000000011111111100011100000000000000110,64'b0000000000000000000000001000000001001111111110000000000010000000,64'b0000000000000000000000000000001100000001100111000000001111000000,64'b0000000000000000000000000100011110011111110000111111011011000000,64'b0000000000000000000000000000010000011111000000000100011111000000,64'b0000000000000000000000000000000100000100000000011111111011000000,64'b0000000000000000000000000000000000001100000000001101111111000000,64'b0000000000000000000000000000011111111110000000001111111111000000,64'b0000000000000000000000000000000000010010000000110011111111100000,64'b0000000000000000000000000000011110000100000011111111111111110000,64'b0000000000000000000000000000010000000000000011111111111101111001,64'b0000000000000000000000000000001000000000001111100111001111111111,64'b0000000000000000000000000000001100001000111111001111110000010000,64'b0000000000000000000000000000000000000111111100001100000001110000,64'b0000000000000000000000000000000000000111110000100111110000000000,64'b0000000000000000000000000000000000001111000011110111101110000000,64'b0000000000000000000000000000000000000010000000000011100000000000,64'b0000000000000000000000000000000000110000000110001010000000000000,64'b0000000000000000000000000000011100111000000001100111111111111111,64'b0000000000000000000000000001111111111000000111111001111111111101,64'b0000000000000000000000001010111111111111111111111110001101001101,64'b0000000000000000000000000111111100001111111100011111100100000000,64'b0000000000000000000000000010110011111111111111111111111111111100,64'b0000000000000000000000001110011100000000110000000111111111110001,64'b0000000000000000000000000011100000011100000000000000000111000001,64'b0000000000000000000000011111111111100011100000000000000111011000,64'b0000000000000000000000000000000000000000000000000000000011111000,64'b0000000000000000000000000000000000000000000000000000000010111100,64'b0000000000000000000000000000000000000000000000000000000001111111,64'b0000000000000000000000000000000000000000000000000000000000111110,64'b0000000000000000000000000000000000000000000000000000000000001111};
assign input_o[39] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000111111111111111111111111100000000000000000000000,64'b0011111111100000000000000111111111111110000000000000000000000000,64'b1011001110000000111111111111111111111100001110010000000000000000,64'b1100111111111111000111111111111111111111100011111111000000000000,64'b0111101111100111000000000000000000000111111110111110000000000000,64'b0011111111111001111111111111111111000000000110000000000000000000,64'b1000001111111000011111111111111111100000001111000000000000000000,64'b0000001110001111111111111111001111111111111111111000000000000000,64'b1000010110000011111111111111111011111111111111111110000000000000,64'b1111111000010000000000001110110111111111111111111100000000000000,64'b1111000001111111111000000010111111100011111011111100000000000000,64'b0000000000000011111100000000011111110001111111100000000000000000,64'b0000000000000000111000000011111011111111111011111000000000000000,64'b0000000000000000011110000001111111111111100000000000000000000000,64'b0000000000000111000011000000000000000000000000000000000000000000,64'b0000000000000000000000000000000110000000000000000000000000000000,64'b0000000000000001000000000000111111000000000000000000000000000000,64'b0000000000000000000000000011111100000000000000000000000000000000,64'b0000000000000000000000000000110000000000000000000000000000000000,64'b0000000000000000000000000100000000000000000000000000000000000000,64'b0000000000000000001010000011100000000000000000000000000000000000,64'b0000000110000100001110000000000000000000000000000000000000000000,64'b0000000110000111001110000000000000000000000000000000000000000000,64'b0000000001111111001110000000000000001000000000000000000000000000,64'b0000000011111111111110000000000000000110000000000000000000000000,64'b0000000000011111000010000000000000000000000000000000000000000000,64'b0000000000000001000010000000000000000000000000000000000000000000,64'b0000000000000010000010000000000000000000000000000000000000000000,64'b0000000000000100000010000000000000000000000000000000000000000000,64'b0000000111111111110000011100000000000000000000000000000000000000,64'b0000001011111101111000001110000000000000000000000000000000000000,64'b0000001110000001111000000000000000000011100000000000000000000000,64'b0000001000000111111000000011000000000000000000000000000000000000,64'b0000001000001111111000000000000000000000000000000000000000000000,64'b0000000000000001111100000001111000000000000000000000000000000000,64'b0000000000000000000000001111111000001000000000000000000000000000,64'b0000000000000000000000001111111000001000000000000000000000000000,64'b0000000000000000000000000000000000001000000000000000000000000000,64'b0000000010111111100000111111111110000000000000000000000000000000,64'b0000000011111111000000111110000000110000000000000000000000000000,64'b0000000001111111000000000000000000111000000000000000000000000000,64'b0000000000000000000000111000000000111000000000000000000000000000,64'b0000000000000000000001111111110011000000000000000000000000000000,64'b0000000000000000000000001110000001000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0011000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000001111111100000000000000000000000000000000,64'b1111110000000000000001111111111111111111111111111110000000000000,64'b0000000000000000000000000111111111001111111111111110000000000000,64'b0000000000000000000000011111110000111111111110000000000000000000,64'b0000000000000000000000011111111111000000111111111110000000000000,64'b0000000000000000000000000000001100001100000011111111100000000000,64'b0000000000000000000000000000000000000111111100000000000000000000,64'b0000000000000000000000000000000000011110011111000000000000000000,64'b0000000001000000000000000000000000000000000001111100000000000000};
assign input_o[40] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000001110000000000000000000000000000000000000000,64'b0000001110000000000000001000000000000000000000000000000000000000,64'b1111111111110000000111000000000000000000000000000000000000000000,64'b1001111111000000001011111100000000000000000000000000000000000000,64'b1111111111110000111111111111000000000000000000000000000000000000,64'b1100000000111001111000000011100000000000000000000000000000000000,64'b0011111100000000000000110000000000000000000000000000000000000000,64'b0111100000000000011111111000000000001111111000000000000000000000,64'b0000000000000000000000000000001111110000000000000000000000000000,64'b0011111111100000000000000001111111111111111100000111111111111000,64'b0011001111000000100000000000000101111100000000001111000011111111,64'b0000000000010111110000000000000111101110000000000000000001111111,64'b0011000000010001010000000000000000110110000000000000000000000000,64'b1111111111111101100000000001010000001111000000000000000000000000,64'b1111000000000000000000000001100000001011100000000000000000000000,64'b1011000000000001111111110000000000000101110000000000000000000000,64'b0000000000000001101111111111111111000011110000000000000000000000,64'b0000000000000000000110000000001111111111111000000000000110000000,64'b0000000000000000000000011111000011100000011000000000000000011111,64'b0000000000000000000000000000010000000000011100000000000000000000,64'b0000000000000000000000000000000000000000010111100000000000000000,64'b0011100000001000000000000000000000000000010000000000000000000000,64'b1111111110100000000000000000000000000000110111000000000000011100,64'b1111111110000000000000000000000000000000110000000000000000000000,64'b1111111100000011100000000000000000000001110000000000000000000000,64'b1111101110100000110000000000000000000001110000000000000000000000,64'b1111111011011000100000000000000000000001110000000000000000000000,64'b1111110111100000000000000000000000000001110000000000000000000000,64'b0001110011111101110000000000000000000001110000000000000000000000,64'b0011001100111111101001000000110000000001110000000000000000000000,64'b1111000111000111111111110001111000000001110000000000000000000000,64'b1100000011100001111111110110111111000001110000000000000000000000,64'b1111000001100000000111101000000011111001110000000000000000000000,64'b1111000110100000000011111111111100110000111000000000000000000000,64'b1111011111110000000000111100100110110100111000000000000000000000,64'b1111000000000000000000111110110110110100011000000000000000000000,64'b1011110000111111000111101111101110111001011100000000000000000000,64'b1011111110100100000100000111100110110001011100000000000000000000,64'b1111111111000001111001100001110110010000011100000000000000000000,64'b0011111100111111111110000011111110010000111111110000000000000000,64'b1110000000011111111111000111101110011000001111111100000000000000,64'b0000000000001111111011000011101110000011111111111110000000000000,64'b0000000000011100000000111111101110000000111111111110000000000000,64'b0000000000000011000000111111000111100000000111111110000000000000,64'b0000000000000000000000000000001001110000000111110000000000000000,64'b0000000000000000000000000000011000011000000000000000000000000000,64'b0000000000000000000000000000001000001100000000000000000000000000,64'b0000000000000000000000000000001100000111000000000000000000000000,64'b0000000000000000000000000000000111110000000000000000000000000000,64'b0000000000000000000000000000000001111100000000000000000000000000,64'b0000000000000000000000000000000000001111000000000000000000000000,64'b0000000000010000000000000000000000000000000000000000000000000000,64'b0000000000000000011111000000000010000000000000000000000000000000,64'b0000000011111111110000000000000010000000000000000000000000000000,64'b0000000000000000000000000000000010000000000000000000000000000000,64'b0000000111111100000000000000000010000000000000000000000000000000,64'b0000000000000000000000000000000010000000000000000000000000000000,64'b0000000000000000000000000000000010000000000000000000000000000000};
assign input_o[41] = {64'b0000000000000000000000000000000000000000000000000010000000000000,64'b0000000000000000000000000000000000000000000111111111000000000000,64'b1110000000000000000000000000000000000000000000000110000000000000,64'b1111110000000000000000000000000000000000000111111100000000000000,64'b1111111000000000000000000000000000001000001111111110011100000000,64'b1111100000000000000000000000000000001000000111111111111110000000,64'b1100000000000000000000000000000000001000000000000000000000000000,64'b1111000000000000000000000000000000001000000000000000000000000000,64'b1000000000000000000000000000000000001000000001111111111111000000,64'b1111010000000000000000000000000000001000000011111111111111110000,64'b0011000000000000000000000000000000001000000000000000000000000000,64'b1110000000000000000000000000000000001000000000111111111111100000,64'b1100000000000000000000000000000000000000000000100001000111100000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000011000000000000000000000000001111111100000001111111111111,64'b0000000000000000000000000000000000010000000000000001110001111111,64'b0011111110000000000000000000000000011111110000000000000000111111,64'b1111111100000000000000000000000000000000000000000000000000000000,64'b1110011100000000000000001111111100000000000000000000000000000111,64'b0001111100000000000000000000001111100000000000000000000000000000,64'b0000011000000000000000011111111111110000000000000000000000000000,64'b0000011000000000000000011111111111100000000000000000000000000001,64'b0110011000000000000000000000000000000000000000000000000000111111,64'b1110011000000000000000000001111111100000000000000000000000111111,64'b1110011000000000000000000001111111100000000000000000000000000000,64'b1111011000000000000000000000000000000000000000000000000000000000,64'b1111011000000000000000000000000000001110000000000000000000000000,64'b0111011000000000000000001100000000011100000000000000000000000000,64'b0011100111000001111000111110000000000000000000000000000000000000,64'b0011100011000000010000110000000000000000000000000000000000000000,64'b0011100011000010010000010000000000000000000000000000000000000000,64'b0011000011000010010000000000000000000000000000000000000000000000,64'b0011000000000010010000000000000000000000000000000000000000000000,64'b0010000000000010010000000000000000000000000000000000000000000000,64'b0000000000000010010000000000000000000000000000000000000000000000,64'b0000000000000010010000000000000000000000000000000000000000000000,64'b0000000000000010011000000000000000001000000000000000000000000000,64'b0001111000000001110000000000000000001000000000000000000000000000,64'b0000000000000000000000000000100000011000000000000000000000000000,64'b0000000000111111110000000000101000011100000000000000000000000000,64'b0000000000111111110000000000000000011100000000000000000000000000,64'b0000000000000000000000000000000011011000000000000000000000000000,64'b0000000000010111000000000000000000001000000000000000000000000000,64'b0000000000111111100000000000000000001000000000000000000000000000,64'b0000000000000000000000000000000000001000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000100000000000100000011111111000000000000000000000000000,64'b0000000000110010000000100000011111111000000000000000000000000000,64'b0000000000110010100111100000000000000000000000000000000000000000,64'b0000000000000000100000000000000000000000000000000000000000000000,64'b0000000000000110100000000000000000000000000000000000000000000000,64'b0000000000000110111100000000000000000000000000000000000000000000,64'b0000000000000110111100000000000000000000000000000000000000000000,64'b0000000000000110000000000000000000000000000000000000000000000000,64'b0000000000000011100000000000000000000000000000000000000000000000,64'b0000000000000011100000000000000000000000000000000000000000000000,64'b0000000000000001100000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[42] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000011111111111111111111111111000000000000000000000,64'b0000000000000000000000010000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000001111000000000001111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000111001100000000000000,64'b0000000000000000000000000000000000000000000000000000000000001100,64'b0000000000000000000000000000000000000000000111000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000111111111111111111111000000000000000000000001111111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000001111111111110000000000000000000000000000001111111,64'b1000000000000000001111111111111110000000000000000000000000001111,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000001111000000000000000000000000000000,64'b0000000000100000000111110000111111100000000000000000000000000000,64'b0000000000100000000000010000111111100000000000111111111111111111,64'b0000000000100000000000000010111111100000000000000000000000000000,64'b0000000000000000000111100011001111111111000000111111010000000000,64'b0000000000100010000000000010011111111111000000011111000111111111,64'b0000000000100000000000000110000011100000000000000000000000000000,64'b0000000000100000000000011110000011001000000000000000000000000001,64'b0000000000100000000000011000000000011100000011110000000000000111,64'b0000000000100000000000100000000000000000000111111100000000000000,64'b0000000000100000000000100000000000000000000000000000000000000111,64'b0000000000100000000000100000000000000000000000000000000000000000,64'b0000000000110000000001100000000000000000000000000000000000000000,64'b0000000000110000000001100000000000000000000000000000000000001111,64'b0000000000110000000001100000000000000000000000000000000000000000,64'b0000000000110000000000010000000000000000000000000000000000000000,64'b0000000000110000000000000000000000000000000000000000000000000000,64'b1100000000010000000000000000000000000000000000001100000000000000,64'b0000000000010000000000000000000000000000001111111111000000000000,64'b0000000000010000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000001111111110000000000000,64'b0000000000010011111000000000000000000000000000000000000000000000,64'b1110000000111110000011000000000000000000000000000000000000000000,64'b1011110000001101000000100111100000000000000000000000000000000000,64'b1001111110000011111110011111100000000000000000000000000000000000,64'b1000000111110001111111000000010000000000000000000000000000000000,64'b0001110001111100000011111111000000000000000000000000001110000000,64'b0000011110111111110000001111111100000000000000000000001100000000,64'b0000000111111111111100000001111100010000000000000000001100000000,64'b0000000011111111001111000000111110011100000000000000011100000001,64'b0000000000011111100001111110000110001100011111111111001000011111,64'b0000000000000111100000111111110010001000111111111111100010011111,64'b0000000000000000000111000111101110000000100000000011100001100001,64'b0000000000000000000011111110001111000000000011111110111010000110,64'b0000000000000000000000001111111111100000000000000101110000010011,64'b0000000000000000000000000110011001000000000000000001111110001101,64'b0000000000000000000000000000011011000000000000000000110110001110,64'b0000000000000000000000000000010000000000000000000000100010010110,64'b0000000000000000000000000000000001000000000000000011100000010111,64'b0000000000000000000000000000010001000000000000000111110000110110,64'b0000000000000000000000000000011001000000000000001111110000111111,64'b0000000000000000000000000000011001000000000000011111110000111110,64'b0000000000000000000000000000011000000000000000001111110010111110,64'b0000000000000000000000000000001000100000000000111111110001111110,64'b0000000000000000001111111111000000100000000001111111110011111110,64'b0000000000000000001111111111000000100000000001001110110011111110,64'b0000000000000001000000100000000111100000000001000110110011111110,64'b0001111100000000011111111111111111100000000000111111110011111110};
assign input_o[43] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000010000000000000000,64'b0000000000000000000000000000000000000000000000010000000000000000,64'b0000000000000000000000000000000000000000000000011000000000000000,64'b0000000000000000000000000000000000000000000000010000000000000000,64'b0000000000000000000000000000000000000000000000010000000000000000,64'b0000000000000000000000000000000000000000000000010000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000111111000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000100000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000011000000000000000000000000000000000000,64'b0000000000000000000000001111110000000000000000000000000000000000,64'b0000000000000000000000010001100000000000000000000000000000000000,64'b0000000000000000000000011111100000000000000000000000000000000000,64'b0000000000000000000000010000000000000000000000000000000000000000,64'b0000000000000000000000010001000000000000000000000000000000000000,64'b0000000000000000000000000001000000000000000000000000000000000000,64'b0000000000000000000000000010000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000011100000000000000000000000000,64'b0000000000000000000000000001000000000000000000000000000000000000,64'b0000000000000000000010001101000000000000000000000000000000000000,64'b0000000000000000000000001101111111111110000000000000000000000000,64'b1100000000000000000000001110000000111110001100000000000000000000,64'b0000000000000000000000000100100111100000011100000000000000000000,64'b0001100000000000000000000100100000000000111100000000000000000000,64'b0000000000000000000000000110111100000000000100000000000000000000,64'b0100000000000000000000000111011000010000000000000000000000000000,64'b1010000000000000000000000001000001100000000000110000000000000000,64'b1010000000000000000000000001111111000000000000000000000000000000,64'b1010000000000000000000000011111111000111100000000000000000000000,64'b1010000000000000000000000111001000101111111000000000000000000000,64'b1010000000000000000000000111010010000001111000000000000000000000,64'b1000000000000000000000000111100001111111111110000000000000000000,64'b0000000000000000000000000001101011111110110000000000000000000000,64'b0000000000000000000000000001110001010110000000000000000000000000,64'b0000000000000000000000000000100000000000000000000000000000000000,64'b0000000000000000000000000000100000000000000000000000000000000000,64'b0000000000000000000000000000100000011110000000000000000000000000,64'b0000000000000000000000000000100100000000000000000000000000000000,64'b0000000000000000000000000000110100100000000000000000000000000000,64'b0000000000000000000000000000001100100000000000000000000000000000,64'b0000000000000000000000000000000000001110000000000000000000000000,64'b0000000000000000000000000000001111000111000000000000000000000000,64'b0000000000000000000000000000000000100000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[44] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000111111110000000000000000000000000000000,64'b0000000000000000000000111111111111000000000000000000000000000000,64'b0000000000000000000000111111111111100000000000000000000000000000,64'b0000000000000000000001110011110111000001110000000000000000000000,64'b0000000000000000000001111100010110000000000000000000000000000000,64'b1000000000000000000011110100011111001111000000000000000000000000,64'b1100000000000000000001110100011111000111000000000000000000000000,64'b1100000000000000000001111100011111000000100011110000000000000000,64'b1100000000000000000011101100010111000000000000000000000000000000,64'b1100000000000000001001111110000111000000000001111100000000001111,64'b0011000000000000000000111111100011000000011111100000111111110011,64'b0001110000000000000000111110100011000000000000000000000000000000,64'b0000000000000000000000001111010011000000000000000000000000000000,64'b0000000000000000000000000111010100000001100000000000000000000000,64'b0000000000000000001111001111111110011111111111111111100000000000,64'b0111111111111110001111111111111111000111111111111100000000000000,64'b0111000000000000000000011111110001111111111110000000000000000000,64'b0000000000000000001111111111110000111111111111111000000000000000,64'b1111111110000000000000011111111000000000111100000000000000000000,64'b1100111111100000000000001111111100000000111000000100000000000000,64'b0000000000000000000000000111111100000000001100000000000000000000,64'b0000000000000000000000000111101100000010000000000000000000000000,64'b0000000000000000000000000101101100100000000000000000000000000000,64'b0000000000000000000000000110111101100000000000000000000000000000,64'b0000000000000000000000000111111100110000000000000000000000000000,64'b0000000000000000000000000111111101100000000000000000000000000000,64'b0000000000000000000000000111001101100000000000000000000000000000,64'b0000000000000000000000000111111101000000000000000000000000000000,64'b0000000000000000000000000011111100111000000000000000000000000000,64'b0000000000000000000000000000000000011000000000000000000000000000,64'b0000000000000000000000000000000000111000000000000000000000000000,64'b0000000000000000000000000000000000011000000000000000000000000000,64'b0000000000000000000000000000000001110000000000000000000000000000,64'b1111101111100000000000000000000000000111111111111111111000000000,64'b1111111111111100000000000000000000011111111111111111111000000000,64'b0000000000000000000000000000000000000000110001111000000000000000,64'b0000000000000000000000000000000000000011111111111111100000000000,64'b0000000000000000000000000000000000000000110000000000000000000000,64'b0000000000000000000000000000001111000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[45] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000111111111111111111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000111111111111111110000011,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000011111111111111111111101111,64'b0000000000000000000000000000000000000001111111111000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000001111110000000000000000010,64'b0000000000000000000000011000000000000001111100000000000000000010,64'b0000000000000000000000000000000000000000001000000000000000000010,64'b0000000000011111000000000000000000000000000000000000000000000010,64'b0000000000101111100000000000000111100000001000000000000000000010,64'b0000000000100011100000000000001111100000000000000000000000000010,64'b0000000000001111000000000000001111100000000000000000000000000010,64'b0000000000000000000000000000000111000000000000000000000000000000,64'b0000001111000000000000000000000111000000000000000000000000000110,64'b0000001111100000000000000000000000000000000000000000000000010011,64'b0000000000000000000000000000000011000000000000001110000000010011,64'b0000000000100000000000000000000111111100000000000000000000010010,64'b0000100000000000000000000000011000111111110000001100000000010110,64'b1001100000000000000000000000000001011111110000000000000000110110,64'b0000001000001000000000000000000001000001110000000000000000110110,64'b0000011100000000000000000000001110000001111000000000000000110110,64'b0000000000000000000000000000001111000001111000000000000000010110,64'b0000000000000000000000000000001111000000111000000000000000010110,64'b0000111111000000000000000000001110000000111000000000000000010110,64'b0001111100111111111111111110011110000000111000000000000000000010,64'b0000011000111111110000000000011100000011100000000000000000000000,64'b0000000000110000001111111111111000000111000000000000000000000000,64'b1111100000110000001111111111111111111111000000000000000000000000,64'b1111100000100000000000000000001111111110000000000000000000000000,64'b1111111110000000000000000000111101111111000000000000000000000000,64'b1111111110000000011100000011111111111100000000000000000000000000,64'b1111101110110000000000000011111111111000000000000000000000000000,64'b1111110111111000000000001111111110000000000000000000000000001111,64'b1111110111111000000000001111111110000000000000000000000000000000,64'b1111100111111000000000001111011100000000000000000000000010000000,64'b1101100110111000000000001111111000000000000000000000001010000000,64'b1111101111110000000000001111110001000000000000000000011010000000,64'b1111001110110000000000011110111001000000000000000000011010000000,64'b1011001101110000000000011110110001000000000000000000001010000000,64'b1011001101100000000000011100010001000000000000000000000010000000,64'b1111001101100000000011111111100000000000000000000000001110000000,64'b1111001101100000000111111101101000000000000000000000000000000000,64'b1110001011100000000011111110000000000000000000000000000000000000,64'b0000000111100000000001111100000000000000000000000000000000000000,64'b0000000000000000000001111000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[46] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000010000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000001000000000000000111100000000000000000000000,64'b1111111111111111111111111110000000000000000000000000000000000000,64'b0000000001111111111110000000000000000000001100000001100000000000,64'b1111111111111111111111111111111111100000000000111111110000000000,64'b0000000000000000111000000000000000000111111111000000000000000000,64'b1111111111111111111111111111111111111111111111111111111100000000,64'b0000000000000000000001110000001110011001111111000000000000000000,64'b0000000000000000000000000001000000010011111111000000000000000000,64'b0000000000000000000000000011111000000001000000000000000000000000,64'b0000000000000000000000111111001100000000000000000000000000000000,64'b0000000000000000000001111111111000000000000000000000000000000000,64'b0000000000000000000011111111111100000000000000000000000000000000,64'b0000000000000000000111111110000000000000000000000000000000000000,64'b0011111111111100111111101110111111110000000000000000000000000000,64'b0000000000000000011100101100111111110000000000000000000000000000,64'b0000000000000000011100111101111111110000000000000000000000000000,64'b0000000000000000011100011111111111100000001100000000000000000000,64'b0000000000000000011101011001101111111000001110000000000000000000,64'b0000000000000000011101000000001111111000111110000000000000000000,64'b0000000000000000011111000111101011101101111110000000000000000000,64'b0000000000000000000111111110011111111111111110000000000000000000,64'b0000000000000000000111111111111111111111111100000000000000000000,64'b0000000000000000000000000011111000010000011100000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000001100000000000000000000000,64'b0000000000000000000000000000000000000000000100000000000000000000,64'b0000000000000000000000000000000010001111111000000000000000000000,64'b0000000000000000000000000000001110011111111000000000000000000000,64'b0000000000000000000000000000011111111111111000000000000000000000,64'b0000000000000000000000000000001110111111111000000000000000000000,64'b0000000000000000000000000000001010111111100100000000000000000000,64'b0000000000000000000000000000011010110011111110000000000000000000,64'b0000000000000000000000000010011111000001111110000000000000000000,64'b0000000000000000000000000001001111111111111111000000000000000000,64'b0000000000000000000000000011101111111000111111000000000000000000,64'b0000000000000000000000000011100010000011111111000000000000000000,64'b0000000000000000000000000000000000000000011111000000000000000000,64'b0000000000000000001111111101100011111100000000000000000000000000,64'b0000000000000000000000000100000000000000000000000000000000000000,64'b0000000000000000000000000010000000000000000000000000000000000000,64'b0000000000000000000000001110000000000000000000000000000000000000,64'b0000000000000000000000001000111100000000000100000000000000000000,64'b0000000000000000000000000001111100000000000000000000000000000000,64'b0000000000000000000000000111001000011111111110000000000000000000,64'b0000000000000000000000001111100000000111111110000000000000000000,64'b0000000000000000000111111011000000000001111100000000000000000000,64'b0000000000000000000001110000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000111111000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[47] = {64'b1100000000000000000000000000000000000010000000000000000000000000,64'b1100000000000000000000000000000000000000100000000000000000000000,64'b1110000000000000000000000000000000000000110001110000100000000000,64'b1110000000000000000000000000000000000000011100110111110000000000,64'b1110000000000000000000000000000000000000011100001101011100000000,64'b1111000000000000000000000000000000000000000100111111111100000000,64'b1111000000000000000000000000000000000000000011111111111100000000,64'b1111000000000000000000000000000000000000000000001111111100000000,64'b1111000000000000000000000000000000000000000000000111111000110000,64'b1111000000000000000000000000000000000000000000001111111000000000,64'b1111000000000000000000000000000000000000000000000100010000000000,64'b1110000001110000000000000000000000000000000000000111111111000010,64'b1110000111111100000000000000000000000000000000000000000000000000,64'b1110000100000000000000000000000000000000000000000000000000000000,64'b1100000011100000000000000000000000000000000000000000000000000001,64'b1110100010000000000000000000000000000000000000000000000000000001,64'b1100000011000000000001110000000000000000000000000000000000000000,64'b1100011110000011000000110000000000000000000000000000000000000000,64'b1100111100011000000000000100000000000000000000000000000000000000,64'b1100000001111111000000001110000000000000000000000000000000000000,64'b1100011111111100000000000011000000000000000000000000000000000000,64'b1100100011111111100000000111000000000000000000000000000000000000,64'b1110001111111011100000000111000000000000000000000000000000000000,64'b1100000011111100111000000111000000000000000000000000000000000000,64'b1100000001110110011110000011000000000000000000000000000000000000,64'b1100011001111110001110000000000000000000000000000000000000000000,64'b1100000000011011110011000000010000000000000000000000000000000000,64'b1100000000001101111101111000011000000000000000000000000000000000,64'b1100001000100100011110011100111100000000000000000000000000000000,64'b1100000000000011010111000110001110000000000000000000000000000000,64'b1100000000001000101101110110000110000000000000000000000000000000,64'b1100000010000000000010110011101110000000000000000000000000000000,64'b1100000010000000000000000100111110000000000000000000000000000000,64'b1100000010000000000000000100001010000000000000000000000000000000,64'b1100001111000001001000000000000111111100000000000000000000000000,64'b1100000011100101101100000000110111111100000000000000000010000000,64'b1100100011111000010011000000100111110110000000000000000000000000,64'b1100100001110011100010000000100111111101000000000000000001000110,64'b1100000001110010101100000000000011011100000000000000000000000000,64'b1100000000111011111100000000000001110011000000000000000000000000,64'b1100000000011111111111100111111100000011001111100000000000000000,64'b1100000000001111111111111110111111000001000000000000000000000000,64'b1100000000000111111111111111111101100001000000000000000000000000,64'b1100000000000000000111111111111111110001100000000000000000000000,64'b1100000000000000000001111111111111010001111000000000000000000000,64'b1100000000000000000000000000000111111010111110000000000000000000,64'b1100000000000000000000000000000001110111111111110010000000000000,64'b1100000000000000000000000000000000111110111111111010000000000000,64'b1100000000000000000000000000000000111111110011011010000000000000,64'b1100000000000000000000000000000000001111111101111110000000000000,64'b1100000000000000000000000000000000000111111111000110000000000000,64'b1100000000000000000000000000000000000001111111111011000000000000,64'b1100000000000000000000000000000000000000111111111000000000000000,64'b1100000000000000000000000000000000000000001111111000000000000000,64'b1100000000000000000000000000000000000000000001110000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000};
assign input_o[48] = {64'b0000000000000100000000000000000000000000000000000000000000000000,64'b0000000000001000000000000000000000000111111111111000000000000000,64'b0000000000001000000000000000000000000000000000001111000000000000,64'b0000000000000000000000000000000000000000000001111000000000000000,64'b0000000000000000000000000000110000000000000111111111010000000011,64'b0000000000000000000000000000000000011000000110011110000000000011,64'b0000000000000000000000000011110000000000000100001010000000111111,64'b0000000000000000000000000011000000000000110000000001111000011110,64'b0000000000000000001110000000000000000000000000000000010000011111,64'b0000000000000001111000000000000001111100000000110000000000011111,64'b0000000000000000000000000000000000000000111101111111111111111110,64'b0000000000000000000000000000000000000011111000000011111100011110,64'b0000000000000000000000000000000000001110000000011111110011111110,64'b0000000000000000000000000000000000011000000000000011111100001100,64'b0000000000000000000000000000001111110000000000011100000000010000,64'b0000000000000000000000000000000111100000011111111111111110011100,64'b0000000000000100000000000000001111111000001111111111000010111110,64'b1111100000000000000011111111111000000000001111111111111111111111,64'b1111110000000000001111111111100111111000011111111111111111111111,64'b0000110000000000011111100000001111110000000000111111000000011100,64'b1111000000000000000000111111111100000000000000000000000000000000,64'b1111000000000011000011111111100000000000000000000000000000000000,64'b0000011100000001000000000000000000000000000000000000000000000000,64'b0010000000000000000000000000000000000000000000000000000000000000,64'b0011100000000000000000000000000000000000000000000000000000000000,64'b1110000000000100000000000000000000000000000000000000000000000000,64'b0000000000000100000000000000000000000000000000000000000000000000,64'b0001111111111100000000000000000000000000000000000000000000000000,64'b0011111111100000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1111111110000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000001000000000000000000000000000011,64'b0000000000000000000000000000000000000000000000000000000000110000,64'b0100000000000000000000000000000000000001100000000000000000000111,64'b1110000000000000000000000000000000000001100000000000000000011111,64'b1111100000000000000000000000000000000010100000000000000001110000,64'b1011110000000000000000000000000000000000100000000000011000000000,64'b1110000000000000000000000000000000000000000000000000011000000000,64'b1110000000000000000000000000000000001100000100000000000000000000,64'b0001100000000000000000000000000000001100000110000000000000000111,64'b0001100000000000000000000000000001001010000110000000000000011111,64'b0000000000000000000000000100000001000000000100000000000011111111,64'b0000000000000000000000001011110001110111111011111111111111110000,64'b0000000000000000000000000000000001100000001001111111111100001110,64'b0000000000000000000000000011110001000000001000001111010001001110,64'b0000000000000000000000000000000001000000001000000011111111100000,64'b0000000000000000000000000000111110000111110000111111111110000000,64'b0000000001111100000110000001111100001111111100000000000000000000,64'b0001111111111100000000000000000000011111100110000000000000000000,64'b0001000111111000000000000000000000000000000100000000000000000000,64'b0000000000000100000000000000000000000011100000000000000000000000,64'b0000000000000100000000000111100000001001100000000000000000000000,64'b0000000011100100100000000111111000011001111000000000000000001010,64'b0000000000000100000000000000000000000000000001111110000000001010,64'b0000000000000100000000000100000011111000000000111000000000001000,64'b0000000000000000000000001100000001001000000000011000000000001000,64'b0000000000000000000000001100001001100000000011111000000000000000,64'b0000000000000000000000000000000000000000000000110000000000110000,64'b0000000000000000000000000010000000000000000000000000000000010000,64'b0000000000000000000000000111000000000000000000000000000000000010,64'b0000000000000000000101111010000000000000000000000000000000000010,64'b0000000000000000000101110000001100000000000000000000000000000000,64'b0000000000000001100011100000000000000000000011000000000000000000};
assign input_o[49] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000111111100000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000011111111111000000000000000000000,64'b0000000000000000000000000001111111111111111111000000000000000000,64'b0000000000000000000000000000111111111111100011000000000000000000,64'b0000000000000000000000111111111111111111111111100000000000000000,64'b0000000000000000000011111100000000000000000001110000000000000000,64'b0000000000000011000000011000000000000000000000111000000000000000,64'b0000000000000000000110111000000000000000000000111000000000000000,64'b0000000000000111100000110000000000000000000000110000000000000000,64'b0000000000000011100000110000000000000000000000110000000000000000,64'b0000000000000111111111100000000000000000000000110000000000000000,64'b0000000000001100000111000000000000000000000000011000000000000000,64'b0000000000011111111110000000000000000000000000011000000000000000,64'b0000000000111100111110000100000000000000000000011000000000000000,64'b0000000000001111111111111000000000000000000001110000000000000000,64'b0000000011110111111111111000000000000000000000011100000000000000,64'b0000000000110001111111111000000000000000000000001100000000000000,64'b0000000000110001111111110000000000000000000000000000000000000000,64'b0000000010000000000010010000000000000000000000001000000000000000,64'b0000000111000000000000010000000000000000000000001000000000000000,64'b0000000110000000000000000000000000000000000000001000000000000000,64'b0000001110000000000101100000000000000000000000000000000000000000,64'b0000001100000000000110110000000000000000000000000000000000000000,64'b0000011000000000000110100000000000000000000000000000000000000000,64'b0000000000000001111111100000000000000000000011011000000000000000,64'b0000000000000011110001100001010000000000000011100000000000000000,64'b0000000111111111111101100001110000000001111100000000000000000000,64'b0000001111111111011111100011010000000001100100000000000000000000,64'b0000000000000001101101000011010000000001000000000000000000000000,64'b0000000000011111111111100010010000000001000000000000000000000000,64'b0000000000000000110000000110010000000001000000000000000000000000,64'b0000000000000000110000000110010000001110000000000000000000000000,64'b0000000000000000011000001101010000001110000000000000000000000000,64'b0000000000000000011110001101010000001100000000000000000000000000,64'b0000000000000000000000001111100000001000000000000000000000000000,64'b0000000000000000100111111011000000000000000000000000000000000000,64'b0000000000000000000001111001000000000000000000000000000000000000,64'b0000000000000000000111111001100000000000000000000000000000000000,64'b0000000000000000000000000000100001000000000000000000000000000000,64'b0000000000000000000000000000010001000000000000000000000000000000,64'b0000000000000000000000000000010001000000000000000000000000000000,64'b0000000000000000000000000000001111000000000000000000000000000000,64'b0000000000000000000000000000001110000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[50] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000111111111,64'b0000000000000000000000000000000000000111111111111111111111111000,64'b0000000000000000000000111111000011111111111111111110011111111111,64'b0000000001100000000011111111111111111011111111111111111111111111,64'b0000000000000111111111100000111111111111111111111111111111110000,64'b0000000011111111111001111111111111111111111111000000000000000000,64'b0001111111111111111111111111111000000000000000000000000000000000,64'b0000111111111111110000000000000000000000000000000000000000000000,64'b0000000000000111100000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000001111000000000000000000000000000000000000000000,64'b0000000000000000001111100000000000000000000000000000000000000000,64'b0000000000000000001001100000000000000000000000000000000000000000,64'b0000000000000000000100111110000000000000000000000000000000000000,64'b0000000000000000001000000011100000000000000000000000000000000000,64'b0000000000000000000111111100110000000000000000000000000000000000,64'b0000000000000000000000000011110000000000000000000000000000000000,64'b0000000000000000000000110001111000000000000000000000000000000000,64'b0000000000000000000001111001011100000000000000000000000000000000,64'b0000000000000000001110000000111100000000000000000000000000000000,64'b0000111110001111100000000000101100000000000000000000000000000000,64'b0000111111111100000000000000101100000000000000000000000000000000,64'b0111111111000000000000000000101100000000000000000000000000000000,64'b1110000000000000000000000000001110000000000000000000000000000000,64'b0000000000000000000001000000010110000000000000000000000100000000,64'b0000000000000000000001000001010110000000000110000000000000000000,64'b0000000000000000000000100001010110000000000000000000000111111111,64'b0000000000000000000000100001010110000000000000000000000111110111,64'b0000000000000000000000100001010110000000000000000000000111110110,64'b0000000000000000000000100001010110000000000000000000000011001110,64'b0000000000000000000000100000000011000000000001111011110001011100,64'b0000000000000000000000100000000011000000000111111011100001101000,64'b0000000000000000000000000001111011100000000001110001000001111110,64'b0000000000000000000000000111000001100000000000110001000001111010,64'b0000000000000000000011111111110001100000000000000000000001111010,64'b0000000000000000000011101111111100111110000000000000000001111010,64'b0000000000000000000011111100111000001100000000000000000001011010,64'b0000000000000000000011011100001100000110000000000000000001000010,64'b0000000000000000000011011100011111010110001000000000000000000000,64'b0000000000000000000111111101100011100011100000000000000000000001,64'b0000000000000000000110111000000000100011111000000000000000000000,64'b0000000000000000000111111000000000111000011111111100000000000000,64'b0000000000000000000001110000000000011000011110000000000000000000,64'b0000000000000000001001000000000000011111001111111110000000000000,64'b0000000000000000011111100000111100011011100000000011111111100000,64'b0000000000001111011011001110001100010111011111111111111000000000,64'b0000111111111111100011000000111100001001100111111100001110000111,64'b1110000000011100000111000000000001110000001000011111111111110000,64'b0000001111111111111001111111111100000000001111111111111100000000,64'b1100000000000000100111111111000000110111110000000000000000000000,64'b0000000000000000011000000011111111111111000000000000000000000000,64'b0000000000001110011111111111000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[51] = {64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000111111111000000000000000000,64'b1111100000000000000000000000000000011111111111000000000000000000,64'b1111110000000000000000000000000000000000000100001111000000000001,64'b1111101111111000000000000000000000000001111111111111000000001111,64'b1111011111111100000000000000000000000010000111111111000000000000,64'b1111111111100000000000000000000011111111000011111111111100000000,64'b1111111111000000000000000011111110000111111111111111000000000000,64'b1111111111000000000111111111111111110011111111111110000000000000,64'b1111111111000000000000000000001000000111111100000000000000000000,64'b1110111111111110011111111111111111111110000000000000000000000000,64'b1111111111111111111000011111110000000000000000000000000000000000,64'b1111111111111100000000011111100000000000000000000000000000000000,64'b1101111000000000000000111111100000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000011,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000011111100000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1111111111111111111111111111100000000000000000000000000000000000,64'b1011111111111111111111111111100000000000000011111111000000000000,64'b0111000000000011111111111110000000000000000000011111100000000000,64'b1011000000000000000000000000000000000000000000000000000000000000,64'b1111000000000001111111111111100000000000000011111111100000000000,64'b1111100000000000000000000000000110000000011111111000000000000000,64'b1111100000000000000011110000000011110000001110000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000001,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000100000000000000000000000000000000000,64'b1111110000000000000000000000111110000000000000000000000000000000,64'b1111110000000000000000000000000111111000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000001100000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000001110000000000000000000000000,64'b1111110000000000000000000000000000011111100000000000000000000000,64'b1111110000000000000000000000000000011110000000000000000000000000,64'b1111110000000000000000000000001111110011000000000000000000000000,64'b1111110000000000000000000000111110000000000000000000000000000000,64'b1111110000000000000000000000111000000000000000000000000000000000,64'b1111110000000000000000000111101000000000000000000000000000000000,64'b1111111000000000000000111000000000000000000000000000000000000000,64'b1111111000000000000011110000000000000000000000000000000000000000,64'b1111111000000000001111000001100000000000000000000000000000000000,64'b1111111000000011111000000000000000000000000000000000000000000000};
assign input_o[52] = {64'b0001011110111100000000000000100000000000000000000000000000000000,64'b0001111111111111110000011111111111111110000000000000000000000000,64'b0000000111111111111111000001111111100001111110000000000000000000,64'b0000000000001111111111110000000011111110011111110100000000000000,64'b0000000000000000111111100000000000000111111101111110000000000000,64'b0000000000000000000000011110000000000000001111111101110000000000,64'b0000000000000000000000111111111000000000000001111111111111111110,64'b0000000000000000000000011111111111100010011100000111111111101111,64'b0000000000000000000000011000100011000000011111100000001111111110,64'b0000000000000000000000001111100011000011111111111111000000001111,64'b0000000000000000000000001110111111111110000011111011111111000000,64'b0000000000000000000000101111111111111111111100011000011111111111,64'b0000000000000000011111110111111111100111111111000011111111111111,64'b0000000000000100111111110011111100111111111111100000000111111111,64'b0000000000001111000111100111111111011111111111110000000000001111,64'b0000000000011110000001111111111111011010000000000000000000000000,64'b0000000000011111110001100000011111111110111111000000000000000000,64'b0000000000001111111111111001100111111110001001000000000000000000,64'b0000000000001111111111100111111111111100011111000000000000000000,64'b0000000000000111111111100001111100001101111111000000000000000000,64'b0000000000000001111000100011110111111111110111000000000000000000,64'b0000000000000000110010000110110011111111100101000000000000000000,64'b0000000000000000010010000000011111111111001101000000000000000000,64'b0000000000000000000100010110001111111001111101000000000000000000,64'b0000000000000000001110000000110111111111111001000110000000000000,64'b0000000000000000000000001100011111111110000001000011000000000000,64'b0000000000000000000000000000101111111111110000000000000000000000,64'b0000000000000000001110000001110111111110001000001000000000000000,64'b0000000000000000001110000000011101001000000000000000010000000010,64'b0000000000000000111100110000011101011000000001000100010000000010,64'b0000000000000000011000001100001111111111100000000111000000000011,64'b0000000000000000001100000000001111011111111000000001110010000110,64'b0000000000000000000110000000001001001111101100000000010001000110,64'b0000000000000000000011000000001001000111111110000000000000111111,64'b0000000000000000000000000000001010000111111101100000000100111011,64'b0000000000000000000010111111101110001100001110100000000011001010,64'b0000000000000000000011101001011100001100000111000000000000011110,64'b0000000000000000000001101011111101111110000011100000000000000110,64'b0000000000000000000000101011111111011100000000111000000001111100,64'b0000000000000000000000110011100101111100000000001111000000111100,64'b0000000000000000000110111111100011111101111000000000000011011100,64'b0000000000000000000010011111111000000110110111100111100001011000,64'b0000000000000000000010001110111101110011000000001111110011011000,64'b0000000000000000000000101101111111000000100000000011100011110000,64'b0000000000000000000000001001011001111100000000010001110011110000,64'b0000000000000000000000000001111000001001001000000000010111110000,64'b1000000000000000000000000000000000000011111111111111111111110000,64'b0000000000000000000000000000000000000000111111011111111111100000,64'b1100000000000000000000000000000000000011111111111111111111100000,64'b1100000000000000000000000000000000000011001110000000000000000000,64'b0011100000000000000000000000000000000001111111111111111110000000,64'b0000000000000000000000000000000000000000111111111111111110000000,64'b1111100011000000000000000000000000000000001001111101101110000010,64'b0000000000100000000000000000000000000000001111111111010110000101,64'b0000001100000000000000000000000000000000001110111011111100000010,64'b0000000001100000000000000000000000000000001101101100011100000011,64'b0000000000011100000011000000000000000000001110011011111100000000,64'b0000000000000000000011110000000000000000000000100111111100000000,64'b0000000000000000000000000000000000000000000000000111111001000000,64'b0000000000000000111111110001100000000000000000000011111001000000,64'b0000000000000000000000000000000000000000000000000011110111000000,64'b0000000000000000000000000011100000000000000000000011110111000000,64'b0000000000000000000000000000010100000000000000000111111111000000,64'b0000000000000000000000000000000000000011000000000111101101100000};
assign input_o[53] = {64'b0001111000000000000000000000000000000000000000000000000000000000,64'b1111010000100000000000000000000000000000000000000000000000000000,64'b1111111110000000000000000000000000000000000000000000000000000000,64'b1111111111111000000000000000000000000000000000000000000000000000,64'b1111111111110000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000111111110000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000111000000000000000000000000000011,64'b0000000000000000000000000000001111100000000000000000000000001111,64'b0000000000000000000000000000001101100000000000000001000000000111,64'b0000000000000000000000000000011101100000000000000000000000000011,64'b0000000000000000000000000011111111100000000000000000000000000001,64'b0000000000000000000000000111111111100100000000000000000000000000,64'b0000000000000000000000001111111111011111000000001100000000011110,64'b0000000000000000001111111111111111111111000000000100000000000011,64'b0000000000111111111111111111111111100111111111111111111100001110,64'b0000000000000111111111111101111111111011001110000001000000000000,64'b0000000000000000000000000000010111111110000000011111100000000000,64'b1111111111111111111111111111111111111111000111110000000000000000,64'b0000000000000010000001111111111110111111011111000000000000000000,64'b0000000000000000000000111111111111101111111100000000000000000000,64'b0000000000000000000000001111111110100011000000000000000000000000,64'b0000000000000000000000000110011101111111000000000000000000000000,64'b0111111111111111111111100000000001110111000000000100000000000000,64'b0000000111000000000000000000000100111111000000000000000000000000,64'b0000000000000000000000000000011110011110000000000000000000000000,64'b0000000000000000000000000000111111000000000000000000000000000000,64'b0000000000000000000000001010100001000000000000000000000000000000,64'b0000000000000000000000000111110001100000000000000000000000000000,64'b0000000000000000000000000111011011000000000000000000000000000000,64'b0000000000000000000000000011101110000000000000000000000000000000,64'b0000000000000000000000000001101110000000000000000000000000000000,64'b0000000000000000011111110001101110001100000000000000000000000000,64'b0001111111111111111111111001111100001100000000000000000000000000,64'b0000111111111111100000000011011100000000000000000000000000000000,64'b0000000000000000001111111001111010000100000000000000000000000000,64'b0000111111111111111111111101110000000000000000000000000000000000,64'b0001100011111111111111110000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[54] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000011110000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1011100000000000000000000000000000000000000000000000000000000000,64'b1001100000000000000000000000000000000000000000000000000000000000,64'b1001100000000000000000000000000000000000000000000000000111111111,64'b0111000000000000000000000000000000000000000000000000001111001111,64'b0000000000000000000000000000000000000000000000000000000111111111,64'b0111110000000000000000000000000000000000000111111100011111111111,64'b0000000000000000000000000000000000000000000100000111110000000000,64'b0000000000000011000000000000000000000001100011111111100000000000,64'b0000000000000000000000000000000000000001111111111111000000000000,64'b0000000000000011111000000000000000000011111101110000000000000000,64'b0000000000000000000000000000000000000000111100000000000000000000,64'b0000000000000000000000000000000000000000111100000000000000000000,64'b0000000000000000000000000000000000001001110000000000000000000000,64'b0000000000000111111000110110000010011111110000000000000000000000,64'b0000000001000000111100110000000010011111100000000000000000000000,64'b0000110011000000000000011111100111011111110000000000000000000000,64'b0000000110000000111100001111111111011111000000000000000000000000,64'b0000111100000001111100010111110111111111000000000000000000000000,64'b0011111000111111100000000011100011101111000000000000000000000000,64'b0010000010111111010001000011100111111110000000000000000000000000,64'b0000000111011110111000000011000011111110000000000000000000000000,64'b0000000011100001100000000011000001111100000000000000000000000000,64'b0000000001111101100000000011001000011000000000000000000000000000,64'b0000000001000100000000000011011000000000000000000000000000000000,64'b0000000000000001100000001110111101111100000000000000000000000000,64'b0000000000000001100000011111000001111110000000000000000000000000,64'b0000000000000000000000011101100001110110000000000000000000000000,64'b0000000000000000000000001101100001111110000000000000000000000000,64'b0000000000000000000000001101100001111110000000000000000000000000,64'b0000000001100000000000011111101001111111000000000000000000000000,64'b0000000000001000000000111111100001111111000000000000000000000000,64'b0000000000000000000000111011100001111111000000000000000000000000,64'b0000000000000000000000001111000001111110000000000000000000000000,64'b0000000000100000000000001111000000011100000000000000000000000000,64'b0000000000111000000000000000000111001110000000000000000000000000,64'b0000000000000000000000000000000111011110000000000000000000000000,64'b0000000000000000000000000000000100000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000111,64'b0000000000000000000000000000000000000000000000000000000011111110,64'b0000000000000000000000000000000000000000000000000000000111111100,64'b0000000000000000000000000000000000000000000000000011111110001111,64'b0000000000000000000000000000000000000000000000011111111011111110,64'b0000000000000000000000000000000000000000000001111111000111110000,64'b0000000000000000000000000000000000000000001111111011111100000000,64'b0000000000000000000000000000000000000001111111101111110000000000};
assign input_o[55] = {64'b1000111011110000000000000000000000000000000000000000000000000000,64'b0111111111100000000000000000000000000000000000000000000000000000,64'b0111000111100000000000000000000000000000000000000000000000000000,64'b1001110111000100000000000000000000000000000000000000000000000000,64'b1010000000000000000000000000000000000000000000000000000000000000,64'b1110011000000000000000000000000000000000000000000000000000000000,64'b0110111100000000000000000000000000000000000000000000000000000000,64'b0011011100000000000000000000000000000000000000000000000000000000,64'b1111011100000000000000000000000001000000000000000000000000000000,64'b1111101111000000000000000000000011110000000000000000000000000000,64'b0001110111000000010000000000000111110000000000000000100110000000,64'b0000111110000000000000000000000110110000000000000000111111000000,64'b0000011110000000001010000000000011110000000000000000111111000000,64'b0000000000000000010110100000000000101111111100000000011111000000,64'b0000000000000000011111110000000000011111111100000000011110000000,64'b0000000000000000010001110000000000000111110000000000000110000000,64'b0000000000000000011111111111000111011111111100000000000000000000,64'b0000000000000000000001111001000011111110001100000000000000000000,64'b0000000000000000000111110000000011111111111100000000000000000000,64'b0000000000000000000000001111110111111111111100010000000000000000,64'b0000000000000000000000000001111111111100000011111000000000000000,64'b0000000000000000000000000000001111111100000001011000000000000000,64'b0000000000000000000000000000000011111000000001111000000000000000,64'b0000000000000000000000001111110001111000000010111100000000000000,64'b0000000000000000000000111111111000011100000001111100000000000000,64'b0000000000000000000000111101001110011101110000000000000000000000,64'b0000000000000000000000110000111111101111111100000000000000000000,64'b0000000000000000000000001111011111111111110110000000000000000000,64'b0000000000000000000000000001111011111111110011110000000000000000,64'b0000000000000000000000011000011110110001111101111100000001111110,64'b0000000000000000000000010000011111101001110000111111111011111111,64'b0000000000000000000000000000000011100010011001111111111110111000,64'b0000000000000000000000000000000001110000011001110100000010111110,64'b0000000000000000000000000000000000100000001110111100000000000000,64'b0000000000000000000000000000000000000000000110000000000001111111,64'b0000000000000000000000000000000001111001110000010000000000000110,64'b0000000000000000000000000000000000000010001110000000000000000000,64'b0000000000000000000000000000000001111110001110000000000000000000,64'b0000000000000000000000000000000001111110001110000000001111111000,64'b0000000000000000000000000000000001111110001110000000000001101100,64'b0000000000000000000000000000000000111011000011000000111110000000,64'b0000000000000000000000000000000000111111000011001000011111100000,64'b0000000000010000000000000000000000111111100001001101101111110000,64'b0000001111111110000000000000000000111011100001001001100000000000,64'b0000000001111111110011111100000000011111100001001000100000000000,64'b0000000111111000000111110011110000000001110000000000011000000000,64'b0000000000001111110111111110001100000000110000111000000000000000,64'b0000000000011111111000011111111000000010110000011110000001111110,64'b0000000000011110111000000011111111101111100000000000000011111100,64'b0000000000001111111000000000000110011111110111000000000000111111,64'b0000000000000011111000000000011100000011110101000000000000111111,64'b0000000000000011110000000001111100000000000111000000000000000000,64'b0000000000000000001111111111111100000001100000000000000000000000,64'b0000000000000000111111111111110100000000111000000000000000000000,64'b0000000000000000111101101111100110011000000000000000000000000000,64'b0000000000000000011011111111110110000000011000000000000000000000,64'b0000000001111111111011111000000110000000000000000000000000000000,64'b0000001111111111110000000000000110000000000000000000000000000000,64'b0000000111100111110100000000000110000000000000000000000000000000,64'b0000011111101101000000000000000111000000000000000000000000000000,64'b0000011111111111000110000111110110000000000000000000000000000000,64'b0000011110111100111111000111110110011110000000000000000000000000,64'b0000001111100100011110000000111110011111000000000000000000000110,64'b0010001111011100001111100000100000011111000000000000000000000000};
assign input_o[56] = {64'b0000000000000000000000000000000000000000000000000000000000010000,64'b0000000000000000000000000000000000000000000000000000000000011111,64'b0000000000000000000000000000000000000000000000000000000101110000,64'b0000000000000000000000000000000000000000000000000000111100110000,64'b0000000000000000000000000000000000000000000000000000001000110000,64'b0000000000000000000000000000000000000000000000000000111100000000,64'b0000000000000000000000000000000000000000000000000000000101000111,64'b0000000000000000000000000000000000000000001111111000111110001111,64'b0000000000000000000000000000000000000000001000011001100000001111,64'b0000000000000000000000000000000000000000011111101110111000000001,64'b0000000000000000000000000000000000000000111111111110011100011111,64'b0000000000000000000000000000000000000011110000000011110110001111,64'b0000000000000000000000000000000000000011100000000011001100000111,64'b0000000000000000000000000000000000000011100000000110010111111111,64'b0000000000000000000000000000000000000111000000000111011100111010,64'b0000000000000000000000000000000000001110100000000011111100111111,64'b0000000000000000000000000000000000001110000000000111100110011010,64'b0000000000000000000000000000000000000111100001111111000010011010,64'b0000000000000000000000000000000000000011110000111100000001110111,64'b0000000000000000000000000000000000000110110001110000000000111111,64'b0000000000000000000000000000000000000110101011110011111100000010,64'b0000000000000000000000000000000000111110010111110111111011011110,64'b0000000000000000000000000000000001111111111111111111111111111111,64'b0000000000000000000000000000000011001111111111000111000110100010,64'b0000000000000000000000000000011110000111000000000001100111011110,64'b0000000000000000000000000000011110000001110000000001111111000001,64'b0000000000000000000000000111111000010000110001000000111101111000,64'b0000000000000000000000001110000000000000010000000000000011111111,64'b0000000000000000000000011100010000000111110000000000000011111011,64'b0000000000000000000000010111100111111111100000000000000000111111,64'b0000000000000000000000001100011111111000000000000000000000011101,64'b0000000000000000000001001011100000000000000000000000000000000101,64'b0000000000000000000000000011000000000000000000000000000000000111,64'b0000000000000000000000111000000000000000000000000000000000001110,64'b0000000000000000000011100000000000000000000000000000011000011011,64'b0000000000000000001100000000000000000000000000000001111010000111,64'b0000000000000011111000010000000000000000000000000001111100000000,64'b0000000000001111101111111100000000000000000000000011110000000000,64'b0000000001111100111111111100000000000000000000000001110000000011,64'b0000000111100011111111111100000000000000000000000111000101000111,64'b0000001111011011111100100000000000000000000000011000000000011110,64'b0000011111111111101000010000000000000000000000000000000000111000,64'b0000001011110000001000010000000000000000000000000000000011111000,64'b0000000110000000011110000000000000000000000010000000000111000011,64'b0000000100000000111000000000000000000000000110000001111110111110,64'b0000000000000000011100000000000000000000101000000101111111110000,64'b0000000000000000011100000000000000000001111000001111110010011100,64'b1111111111111111111111111111111111111111111111111110010000001100,64'b1111111111111111111111111111111111111111111111111111100000001111,64'b1111111111111111111111111111111111111111111111111111000001111100,64'b1111111111111111111111111111111110111111011111101111000001100000,64'b1111111111110011111111101111111111111111111011111111000111100000,64'b1111110111111111111110111111111111111111111111011111000111110000,64'b1110111111111011111111011111111110111111111111111011100110010000,64'b1111111111111111111111111111111111111111111111100001111110110000,64'b0000000000000011000010011001000000000011011000000000111110110000,64'b1000000000000011000000000111000000000001101110000000000001000001,64'b0000000000000110000000000011000000000001110110000000000001100000,64'b0000000000000111000000000011000000000000110111000000000001100000,64'b0000000000000111000000000110000000000000100101100000000001100000,64'b0000000000001110000000000110000000000000001001100000000011000000,64'b0000000000001100000000001110000000000000001100010000000001000000,64'b0000000000001100001000101100000000000000000100001000000001000000,64'b0000000000001100001000111100000000000000000100001000000001010000};
assign input_o[57] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000001111110000000000000,64'b0000000000000000000000000000000000000000011111111110000000000000,64'b0000000000000000000000000000000000000011111110000011111100000000,64'b0000000000000000000000000000000000000000000011010001111111111111,64'b0000000000000000010000011111110000000000000000001100000001111111,64'b0000000000000000011100000000100000000000000000000000001000000000,64'b0000000000000000001111100000100000000000000000000000000000000011,64'b0000000000000000000001100001100000000000000000000000000000000000,64'b0000000000000000011001111111111111000000000000000000000000000000,64'b0000000000000000010000000000000000000000000000000000000000000000,64'b0000000000000000000111001111111110000000000000000000000000000000,64'b0000000000001100110001000000000000000000000000000000000000000000,64'b0000000000000000000000111111100000000000000000000000000000000000,64'b0000000000000000000011000011100000000000000000000000000000000101,64'b0000000100000000000001001000000000000000000000000000000000000011,64'b0000000000000000000000111111100000000000000000000000000000000111,64'b0000000000000000000010000111100000000000000000000000000000000111,64'b0000000000000000000010000000000000000000000000000000000001111111,64'b0000000000000000000000000000000000000000000000000000000000011101,64'b0000000000000000000000100100000000000000000000000000001100000110,64'b0000000000000000000001101110000000000000000000000000000000000101,64'b0000000000000000000001001000000000000000011100000000000000000011,64'b0000000000000000000000000011100000000000000011000000000000000000,64'b0000000000000000000000000000000000000000011110000000000000000000,64'b0000000000000100111000001001000000000000001111000000000000000000,64'b0000000000001111111000001101000000000000110000000000000000000000,64'b0000000110001111011010001110000000000110110000000000000000000000,64'b0111111111110000000111000111100000000000011100000000000000000000,64'b1111111100000000001111111111100000000000111110000000000000000000,64'b1000000000000011111011100011111111100000011110000000000000000000,64'b1100000000000111111000001111110100001111111111000000000000000000,64'b1100000000000111001111001111111000000111111111000000000000000000,64'b1110000000000111001110000000111100011011111110110000000000000000,64'b1110000000000011100110000000111000001100110111111000000000000000,64'b1100000000000001100110000000001101001100111000011000000000000000,64'b0011000000000000110011000000001110100111110000000000000000000000,64'b1111000000000000111011100000000111000110001100000000000000000000,64'b1111000000000000111001111111111101100000000001110000000000000000,64'b0011100000000000011110000000001111000000000011111000000000000000,64'b1111100000000000000110000000000000000001000111100000000000000000,64'b1101100000000000000111111000000000110001000110000000000000000000,64'b0001100000000000000110111100001111110000000111001110000000000000,64'b1111100000000000000111110111111111100000000111110000000000000000,64'b0111110000000000000011111001111111111100000111111110000000000000,64'b0111111100000000000001100000111001001101100010001110000000000000,64'b1110111100000000000001111111100000001010001011111100000000000000,64'b1111111110000000000000111001100000000111000100001100000000000000,64'b1111111110000000000000001111000000000001111111110000000000000000,64'b0011101110000000000000000000001000000000111100000000000000000000,64'b0011111111110000000000001111111000000000111111111100000000000000,64'b1001111011110000000000000111111100000000000000000000000000000000,64'b1100111101111000000000000011111111000001100000000000000000000000,64'b1100011111111000000000000010110110111011000000000000000000000000,64'b1100011110111100000000000000110111111111100000000000000000000000,64'b1111000111001100000000000000111111111100000000000000000000000000,64'b0111000011001100000000000000111111011111110000000000000000000000,64'b0111100011111100000000000000011111111111110000000000000000000000,64'b0011100001111001100000000000011111000000000000000000000000000000};
assign input_o[58] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000011111100000000000000000000000000000,64'b0000000000000000000000000001111111110000000000000000000000000000,64'b0000000000000000000000000111110011111000000000000000000000000000,64'b0000000000000000000000000111111111111100000000000000000000000000,64'b0000000000000000000000000111110000111100000000000000000000000000,64'b0000001111000000000000000011110000011100000000000000000000000000,64'b1111111111111100000000000001111110011100000000000000000000000000,64'b1111110000001111000000000000111111111000000000000000000000000000,64'b0011110000001111110000000000010000110000000000000000000000000000,64'b0000000000000100010000000000000000000000000000000000000000000000,64'b0000000000000101000000000000000000000000000000000000000000000000,64'b0000000000000111000000000000000000000000000000000000000000000000,64'b0000000000000011100000000000000000000000000000000000000000000000,64'b0000000000000011000000000000000000000000000000010000000000000000,64'b0000000000000110001111000000000000000000000111111000000000000000,64'b0000000000001110001111000000000000000000001000000000000000000000,64'b0000000011111110011011000000000000000000011110100000000000000000,64'b0000000011111100111110000000000000000000011110000000000000000000,64'b0000001111111100110110000000000000000000011011000000000000000000,64'b1111111111111000110110000000000000000000011011000000000000000000,64'b0011111111110000110110000000000000000000011010000000000000000000,64'b0000000000000000110100000000000000000000011010000000000000001111,64'b0000000000000001100100000000000000000000000111000000000001111111,64'b0000000000000001100100000000000000000000000111100000000011110111,64'b0000000000000001100100000000000000000000011000000000000011111111,64'b0000000000000001100100000000000000000001111111110000000001110000,64'b0000000000000000000110000000000000000001111011111000000000110000,64'b0000000000000000001111000000000000000000111111111111111000000111,64'b0000000000000000011111000000000000000000010000111011111100000000,64'b0000000000000001111111100000000000000000000000001111101110000000,64'b0000000000000001110110100000000000000000000000000001111100000000,64'b0000000000000001111110000000000000000000000000000000000000000000,64'b0000000000000000111100000000000000000000000000000000110000000000,64'b0000000000000000010110000000000000000000000000000001011000000000,64'b0000000000000000000010000000000000000000000000000001011000000000,64'b0000000000000001100010000000000000000000000000000001010000000000,64'b0000000000000001100110000000000000000000000000000001010000000000,64'b0000000000000001100010000000000000000000000000000000000000000000,64'b0000000000000001001010000000000000000000000000000000000000001000,64'b0000000000000101011000000000000000000000000000000000000000000000,64'b0000000000000111011000000000000000000000000000000000000000000000,64'b0000000000000111011000000000001000000000000000000000000000000000,64'b0000000000000111011000000000000000000000000000000000000000000000,64'b0000000000000100011000000000000000000000000000000000000000000000,64'b0000000000000100111000000000000000000000000000000000000000000000,64'b0000000000001100110000000000010000000000000000000000000000000000,64'b0000000000001100110000000000010000000000000000000000000000000000,64'b0000000000001100000000000000000000000000000000000000000000000000,64'b0000000000011111000000000000000000000000000000000000000000000000,64'b0000000000011111000000000000000000000000000000000000000000000000,64'b0000000000011111000000000000000000000000000000000000000000000000,64'b0000000000011011000000000000000000000000000000000000000000000000,64'b0000000001111111000000000000000000000000000000000000000000000000};
assign input_o[59] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000001111111111111111111111111,64'b0000000000000000000000000000000111100000011111111111000000000000,64'b0000000000000000000000000000000011000000000000000000111111111111,64'b0000000000000000000000000000000000000000000111111111111111111111,64'b0000000000000000000000000000000000000011111111111111111111111111,64'b0000000000000000000000000001000000011111111111111111001111111111,64'b0000000000000000000000000000000011110000111111111111111111111111,64'b0001111101110000000000000000000000001111111111111111111111111100,64'b0011111111110000000000000000000000001111111110000000000000000000,64'b0000000011110000000000000000000011111111110000000000000000001000,64'b0011111111110000000000000000000000000000000000000000000000000000,64'b0000111111000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000111,64'b1000000000000000000000000000000000000000000000000000000001111111,64'b0000000000000000000000000000000000000000000011111111111111111111,64'b1000000000000001000000000000000000000111111111111111111111111011,64'b0000000001111111111000000000000011111111111111111111111100000001,64'b0000011111111111110000000000001111111111100000011111111111000000,64'b0000001111111000000000000000001111111010111111100000000000000000,64'b0000000111111000000000000000000000111111000000000000000000000000,64'b0000000011100000000000000000000000111111000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000001111000000000000000000000000,64'b0000000000000000000000000000000000001111000000000000000000000000,64'b0000000000000000000000000001111111111000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000111111100,64'b0000000000000000000000000000000000000000000000000001111111000000,64'b0000000000000000000000000000000000000000000001111111110000000000,64'b0000000000000000000000000000000000000000000011111110000000000000,64'b0000000000000000000000000001111111111111111111000000000000000000,64'b1111100000000000000000000000101111100000011000000000000000000000,64'b0000000000000000000000001111111100000000000000000000000000000000,64'b0000000011110000000111111111000100000000000000000000000000000000,64'b1111111110000000111111100000000100000000000000000000000000000000,64'b1111100111111111111000000000000000000000000000000000000000000000,64'b1111111111111111000000000000111100000000000000000000000000000000,64'b1111111111111110000000000000000000000000000000000000000000000000,64'b1111000000000000000000110000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000001100000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[60] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000010000000000000000000000000000000000000000000000000000,64'b0000000000010000000000000000000000000000000000000000000000000000,64'b0000000000010000000000000000000000000000000000000000000000000000,64'b0000000000010000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000010000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000011100000000000000000000000000000000000000000000000000001100,64'b0000011111000000000000000011111111110000011111111000000000000000,64'b0000011011100000000000000011111110000000001111110000000000000000,64'b0000001001100000000000000111001000000000000001110000000000011111,64'b0000000011000000000000000011100000000000000000011000000000000000,64'b1111110000000111100000000001000000000000001111100000000000000000,64'b1111000000001111110000000000000000011100000011110000000000000000,64'b0110001110000010100000000000000000011100000000000001000000000000,64'b1011101110010010000000000000000000011100000000000011111100000000,64'b1111100000010000100000000000000000011100011111000000000000000000,64'b1011100000011100100000000000000000111100110110000000000000000000,64'b1011100000001100100000000000000000111100110000000000000000000000,64'b1011100000011100110000000000000000111100010000000000000000000000,64'b0011000000001100111000000000000000111100000000000000000000000000,64'b0010000000001100111000000000000000111100000000000000000000000000,64'b0010000000001100110000000000000000111100000000000000000000000000,64'b0010000000000011100000000000001001111100010000000000111000000000,64'b1011111111111111100000000000000000111100000000000001111100000000,64'b1100111111111111100000000000001000111100000010011111111000000000,64'b1111111100111110000000000001000000011100000011111000001000000000,64'b0001111111111111000000000001000110011100000011000000011000000000,64'b0000011111111100000000000001000011011100000011110000011000000000,64'b0000000001110000000000000001000010001100000011100000011000000000,64'b0000000000000000000000000001000010001100000001100000011000000000,64'b1000000101101000000000000001000010011000000000100100001110000000,64'b0000000101100010000000000001000000011000000000100100000110000000,64'b0010011101110010000000000001000000011000000000100001000010000000,64'b0011011000110011000000000000100000011000000000100000000010000000,64'b1011011000110011000000000000111010011000000000000000000000000000,64'b1011111000110011000000000000001110011000000000000000000000000000,64'b1011011000110011000000000000000110011000000000000000000000000000,64'b1010011000010010000000000000000010010000000000001000000000000000,64'b1100000000000000000000000000000000110000000000000000000000000000,64'b0000110000000000000000000000000000000000000000000000000000000000,64'b0001100001000011111000000000000000000000000000000000010000000000,64'b0000000001000000000000000000000000000001111110000000000000000000,64'b0000000111111000000000000000000000000001111000000000000000000000,64'b0000001101111011100000000000000011110000000000000000000000000000,64'b0000000001011000000000000000011110000001111110000000000000000000,64'b0000000000110000000000000111111000000000000000000000000000000000,64'b0000011111100000011100000111100000010000000000000000000000000000,64'b0000011110000000011111000111111111000000000000000000000000000000,64'b1000000000111000000000000111110000000000000000000000000000000000,64'b0000000111111100001111110000000000000000000000000000000000000000,64'b0000000001000000001111100000000000000000000000000000000000000000,64'b1111111111111111000000000000000000000000000000000000000000000000,64'b0011111111111000000000000000000000000000000000000000000000000000,64'b1111111111000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[61] = {64'b0000100000000000000000000000000000000000000000000000000000000000,64'b0000110000000000000000000000000000000000000000000000000000000000,64'b0000111000000000000000000000000000000000000000000000000000000000,64'b0000111000000000000000000000000000000000000000000000000000000000,64'b0000010000000000000000000000000000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000000000000000000000000,64'b1111111100000000000000001100000000000000000110000000000000000000,64'b0000001110001111111000000000000000000000000000000000000000000000,64'b0000000000000011111100000000000100000000000000000100000000010000,64'b0000000000000000000000000000000000000000000000000100011000000000,64'b0001110000000011111000000000001100000000000000000000111000000000,64'b0000010000000001111110010010011110000000000000000010111000000000,64'b0000000000000000000000000000000001111111100000000011111000000000,64'b0000000000000000000000000000000000000000111110000011011000000000,64'b0000000000100000000000000000000000000000000010000011010000000000,64'b0000000000110000000000000110000000000000000000000000100000000000,64'b0000001110111000000000000111111100000000000000000010100000000000,64'b0000000111100000000000000000111111110000001111111111110000001110,64'b0000000000000111100000000111111111101111000000000011000000000000,64'b0000000000000001111100000000011111110011000000000011111100100000,64'b0000000000000000000111111100011111111100000010000111111110000000,64'b0000000000001110000000000000001111111111001100000011111111000000,64'b0000000000000000000000000000101100000000001111100011111111000000,64'b0000000000000000001111111111000000000000001111110011111111000000,64'b0000000000000000011111111100000000000000000011111111110111000000,64'b0000000000000000000000000000000000000000000011100100011110000000,64'b0000000000000000000000000000000000000011110010000111001100000000,64'b0000000000000000000000000000000000000011111110000011111000000000,64'b0000000000000000000000000000000000000000011110000011011000000010,64'b0000000000000000000000000000000000111111111001110011111100000010,64'b0000000000000000000000000000000000000000000001000011111100111110,64'b0000000000000000000000000000001111111111000110000011111000000000,64'b0000000000000000000000000000001111111111111110000011111000000000,64'b0000000000000000000000000000011111111111110111010000111000000000,64'b1000000000000000000000000000111111100111110001111111111000000000,64'b0000000000000000000000000000011111111111000001111011111000000000,64'b0000000000000000000100000000011111111111000001111110110000000000,64'b1000000000000000000000000000000111111111100001111111110000000000,64'b1100000000000000000000000000110000001111100001111111111110000000,64'b1100000000000000000000000011111000000011000011111111111111000000,64'b1000010000000111000000000011111100000000000011111111100111000000,64'b0000010100000011100000000011111111101000000010011011100000000000,64'b0000000000000000000000000011111101101000000000011111100000000000,64'b0000000111100000000000000001100101101000000000011111100000001111,64'b0000001111100000000000000000100001111000000000011101100000111111,64'b1000011111100000000000000000000010111000000000001110100000011111,64'b1110011110011111000000000000000011000000000111111111111111111001,64'b1110010100001001111000000000000000000000011110011100111111100111,64'b1110000100000001111000000000000000000000000001111111111111111111,64'b1110001111111111011110000000000000000000001110011111111111111111,64'b1111111111110001111110001000000000000000000000000011111111110000,64'b1111110000000100110110001100000000000000000001000000000000000000,64'b1000000000001111111110011111111100000000001000000000000000000000,64'b0000000000001111000000011111111111000000000000000000000000000000,64'b0000000000000000000000011011110001111000000000000000000000000000,64'b0000000000000000000000011110000011111100000000000000000000000000,64'b0000000000000000000000001111100111111111000000000000000000000000,64'b0000000000000000000000001111111111111111111000000000000000000000,64'b0000000000000000000000000011111111111101111100000000000000000000,64'b0000000000000000000000000000000001111111111111100000000000000000,64'b0000000000000000000000000000000000011111111111111100000000000000,64'b0000000000000000000000000000000000011111111011111110000000000000,64'b0000000000000000000000000000000000001111111111111111110000000000,64'b0000000000000000000000000000000000000001111111110111111000000000};
assign input_o[62] = {64'b0000000000000000000000000000000000000000000000000100000000000000,64'b0000000000000000000000000000010111100011111100010110000000000000,64'b0000000000000000001000000000011111111000000011000110000000000010,64'b0000000000000000000000000000011111111110000001000100000000000010,64'b0000000000000000000000000000011111011100000000111000000000000010,64'b0000000000000000000000000000011111111100000000000000000000000010,64'b0000000000000000000000000000011101011100000000000000000000000010,64'b0000000000000000000000000000011001011100000000000000000000000010,64'b0000000000000000000000000000000110011000000000000000000000000000,64'b0000000000000000000000000000000110110000000000000000000000000000,64'b0000000000000000000000000000000010010000000000000001111111000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000011100011,64'b0000000000000000000000000000000000100000000000000000000111111111,64'b0000000000000000000000000000000000000000000000000000011101111011,64'b0000000000000000000000000000011110000000000000000000000111111111,64'b0000000000000000000000000000111111100000000000000000011111111111,64'b0000000000000000000000000000111011100000000000000000000000011110,64'b0000000000000000000000000000111001100000000000000000000000000010,64'b0000000000000000000000000000101001100000000000000000000000000010,64'b0000000000000000000000000001111111111111000000000000000000000110,64'b0000000000000000000000000011111101111111110000000000000010000010,64'b0000000000000000000000001111110001111111111000000000000000000010,64'b0000000000000000000000001111100000011101111100000000000000000000,64'b0000000000000000000000011110000000001110011100000000111110000000,64'b0000000000000000000000111000000000000111111100000011111111000000,64'b0000000000000000000000110000000000000111111110001111111111000000,64'b0000000000000000000000100000000000000011111110011110001111000000,64'b0000000000000000000000100000000000000111110110011100001111000000,64'b0000000000000000000001100000000000001111111010011001001111000000,64'b0000000000000000000001100000000000000011111010010000011111000000,64'b0000000000000000000001100011000000000000001110011111111100001100,64'b0000000000000000000001111111100001000000011111000011111110000000,64'b0000000000000000000001100101111111111111111111100000000000000000,64'b0000000000000000000001101100111100111111111111000000000011111000,64'b0000000000000000000000111100111110000011111111100000001111111100,64'b0000000000000000000000111111111110000111111111000000011111111000,64'b0000000000000000000000011111111101111111111000000000000000000000,64'b0000000000000000000000000000011101111111100000000001011111111000,64'b0000000000000000000000000000011100001111100000000001111111111100,64'b0000000000000000000000000000011110001011100000000000110111111100,64'b0000000000000000000000000000011100001011100000000000110101011000,64'b0000000000000000000000000000001110001001100000000000110101111000,64'b0000000000000000000000000000001111000101100000000000110101111000,64'b0000000000000000000000000000001111000011100000000000110101111000,64'b0000000000000000000000000000001101001111100000000000110101111100,64'b0000000000000000000000000000110010001111110000000000110010011100,64'b0000000000000000000000000000000000111111110000000011111111001101,64'b0000000000000000000000000000000000011111110000000000000010011000,64'b0000000000000000000000000000000000000111110000000001111111111111,64'b0000000000000000000000000000000000000011111111110000000110000111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[63] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000001000,64'b0000000000000000000000000000000000000000000000000000000000001110,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000001111,64'b0000000000000000000000000000000000000000000000000000000000001111,64'b0000000000000000000000000000000100000000000000000000000011111100,64'b0000000000000000000000000000000100000000000000000000000000000000,64'b0000000000000000000000000000000100000000000000000000000000000000,64'b0000000000000000000000000000000100000000000000000000000000000000,64'b0000000000000000000000000000000100000000000000000000001100000000,64'b0000000000000000000000000000000100000000000000000000011100000000,64'b0010100000000000000000000000000100000000000000000000001100000000,64'b1001100000000000000000000000000100000000000000000000001100000000,64'b1101100000000000000000000000000000000000000000000000011100000011,64'b1101100000001001100000000000000000000000000000000000011000000011,64'b1101100000001101110000011111000000000000000000000000001100000000,64'b1101110000001101110001000001100000000000000000000000001100000000,64'b1101110000001101110000000001100100000000000000000000001100000000,64'b1001110000001101110000000000000100000000000000000000001100000000,64'b1111110000001100110000000000000100000000000000000000001100001000,64'b1011100000001100110000000000000000000000000000000000001100001001,64'b0001100000000000010000000000000001000000000000000000001100001000,64'b0001100000000000010000000000000001000000000000000000001100001000,64'b1111110000000000010000000000000001100000000000000001101110000111,64'b0111110000000000010000000000000111110000000000000001101110001111,64'b0111100000000000000000000000000110110000010000000001101110000000,64'b1111000000000000000000000000001111100000000000000001101111000000,64'b1110000000000001110000000000011101100000000000000001111111000011,64'b0000000000000001111100000000000010110000000000000001110111000011,64'b0000000000000000000000000011111000110000000000000000111111001000,64'b0000000000000000000000000011111100000000000011000000101100000000,64'b0000000000000000000000000011100111100000010111000001100100000011,64'b0000000000000000000000000001111011100000011111000000100110000111,64'b0000000000000000000000000000111111001000001111001111000110000000,64'b0000000000000000000000000000100001000000001110001111110010000000,64'b0000000111111111110011011100100110000000001110111111111011111000,64'b0000000000111111100000011110111111000000000000110000010001111111,64'b0000011111111000000000011100111111000000000000100000000000000011,64'b0000000001111000000011111111111111000000000000000000111111000000,64'b0000000000000000000000001100111111000000000000000111111111000000,64'b0000000000000000000000000000011110000000000000001111111110000110,64'b0000000000000000000000000000011111000000000000000001000000000111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[64] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000001111111110000000000000000000000,64'b0000000000000000000000000000011111111111111000000000000000000000,64'b0010000000000000000000000000000000011111111000000000000000000000,64'b0100000000000000000000000000000000000000011000000000000000000000,64'b0000000000000000000000000000000001111111111000000000000000000001,64'b0000000000000000000000000000000000000011000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000111100,64'b0000000000000000000000010000000000000000000000000000000000000100,64'b0000000000000000000000000000000000000000000000000000000111111100,64'b0000000000000000000000000000000000000000000000000000000011111111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000011111101111111111111111111000000000000000000000,64'b0000000000000000001111111111111111111111110000000000000000000000,64'b0000000000000000000011111111111111111111111000000000000000000000,64'b0000000000000000000000111111111111111111111000000000000000000000,64'b0000000000000000000011111111111111111111111000000000000011111111,64'b0000000000000001000011111100000000000001110000000000000001111111,64'b0000000000000001001100000000001111110000000000000000000100000000,64'b0000000000000001000000000000111111110000000000000000000100000000,64'b0000000000000000010000000011111111110000000000000000000100000000,64'b0011000000000000000000000000000000010000000100000000000011100000,64'b0011111110000000000000000000011111110000000000000000000011111100,64'b0011110000000011000000000000000000000000000000000000000000110011,64'b1100000000000000000000000000000000000000000000000000000000110011,64'b0000000111111111000000000000000000000000000000000000000000100000,64'b0001111111110000000000000000000000000000000000000000000000000000,64'b0011111111111111100000000000000000000000000000000000000000000000,64'b0001111111111001000000000000000000000000000000000000000000000000,64'b1111111111111111111111111111111000011100000000000000000000000000,64'b0000000000000000000000000001111000001100000000000000000000000000,64'b0010000000001111111111000000111000001100000000000000000000000010,64'b0000000000000001111111000000111000001100000000000000000000000110,64'b0001110000000001111111100000111000001100000000000000000000000011,64'b0000000000000001100111100000101000001100000000000000000000000001,64'b0000000000000111011011000000001000001100000000000000000000000001,64'b0000000000011111100111100000000000000100000000000000000000000000,64'b0000001110011111111111100000110000000100000000000000000000000000,64'b0000000000001111111111111100110000000000000000000000000000000000,64'b0000000000001111111111000000110000000000000000000000000000000000,64'b0000000000000111111100000000110000000100000000000000000000000000,64'b1111110000110000000000000000110000000000000000000000000000000000,64'b1111100000111000000000000000110000000000000000000000000000000000,64'b1111100000111000000000000000110000000000000000000000000000000000,64'b1111100011111101000000000000011000000000000000000000000000000000,64'b0010000000100100000000000000001110001111111111111100000000000000,64'b1010011100000000000000000000000111111111111111111111000000000000,64'b0000011000100000000000000000000000111111111111110000000000000000,64'b0001111000100100000000000000000000011111111111111111000000000000,64'b0000111000100000000000000000000000000010000111110000000000000000,64'b0000011000100000000000000000000000000000000000000000000000000000,64'b0000011100000000000000000000000000000000000000000000000000000000,64'b0000011000000000011111100000100000000000000000000000000000000000,64'b0000000000000001101000011111110000000000000000000000000000000000,64'b0000000000000001100000000000110000000000000000000000000000000000,64'b0000000001100000111111111111100000000000000000000000000000000000,64'b0000000011110000011111111111100000000000000000000000000000000000,64'b0001111111111100000000000000000000000000000000000000000000000000,64'b0111111111111100000000000000000000000000000000000000000000000000,64'b0011111111110001110000000000000000000000000000000000000000000000,64'b1111111111111100000000000000000000000000000000000000000000000000,64'b1111111111111111000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[65] = {64'b0000000000000000000111110011111011110011000000000011000000000000,64'b0000000000000000000111100001111001110011111000111111000000000000,64'b0000000000000000000001000000111001110011111000111111100011100000,64'b0000000000000000000000000000011001110010111111111111000010100000,64'b0000000000000000000000000111100110110001111111111111111111000011,64'b0000000000000000000000000111111000000000000000000001111111100110,64'b0000000000000000010000011111111000000000000000000000000000000000,64'b0000000000000000010000000000000000000000000000000111111111111110,64'b0000000000000000010000000000100000000000000000000001111111111110,64'b0000000000000000010000000011111100000000000000001111111111111110,64'b0000000000000000010000001111111111000000000000000001111111111110,64'b0000000000000000010000011111111111000000000000000000000000011100,64'b0000000000000000000000111011110111100000000000000011111110000111,64'b0000000000000000000000111111110111000000000000000000001100000000,64'b0000000000000000000000010111111111000000000000000000000000000000,64'b0000000000000000000000001111111111000000000000000000001000000000,64'b0000000000000000000000000011111100000000000000000000000000000000,64'b0000000000000000000000000000011111111000000000000001111111110000,64'b0000000000000000000000001001111111111100000000000011111111111000,64'b0000000000000000000000001000011100110000000000000011001111111000,64'b0000000000000000000000000001111111111100000000000011100111110000,64'b0000000000000000000000000000000010000000000000000011000011110100,64'b0000000000000000000000000000000000000000000000000011011011110000,64'b0000000000000000000000000001011111111110000000000011011011100000,64'b0000000000000000000000000111111111111110000000000001111111100000,64'b0000000000000000000000000001111000111100000000000000111111000000,64'b0000000000000000000000001000000000001100000000000000000000100000,64'b0000000000000000000000000000000001110000000000000000001111100000,64'b0000000000000000000000001000000100000011000000000001011111100000,64'b0000000000000000000000011111111111111111100000000001011111100000,64'b0000000000000000000000000111111110000001100000000000001011100000,64'b0000000000000000010000100011111111000000011000000000001110000000,64'b0000000000000000010011111100011110000011111000000000000110000000,64'b0000000000000000010111111100000000100010011000000000000000000000,64'b0000000000000000011111111111110000100011101000000001000000000000,64'b0000000000000000011001110111111001111010110000000011000000000000,64'b0000000000000000010111111000011100111010000000000001111100000000,64'b0000000000000000011111111111101000011111000000000000111100000000,64'b0000000000000000000111111111101000001110000000000000000000000000,64'b0000000000000000000000000000001000000000000000000000111000000000,64'b0000000000000000000000000000011000000000000000000000000000000000,64'b0000000000000000000000000001011000100000000000000000000000000000,64'b0000000000000000000000000001011000100000000000000000000000000000,64'b0000000000000000000000000001011000000000000000000000000000000000,64'b0000000000000000000000000000011000000000000000000100111111111100,64'b0000000000000000000000000000011000000000000000000111111111111110,64'b0000000000000000000000000000011000000000000000000011111111101000,64'b0000000000000000000000000000100000000000000000000000111111111110,64'b0000000000000000000000000000001111111101111000001111111111111100,64'b0000000000000000000000000000001111111111101000000111111111111110,64'b0000000000000000000000000000000100000000000000000111111111111010,64'b0000000000000000000000000000111111111100000000000111111111111110,64'b0000000000000000000000000000000000000000000000000000111100000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[66] = {64'b1110000000000000000000000000000000000000110000000000000000000000,64'b1110000000000000000100000000000000000000110000000000000000000000,64'b1110000000000000000100000000000000000000010000000000000000000000,64'b1110000000000000000100000000000000000000000000000000000000000000,64'b1110000000000000000011000000000000000000001100000000000000000000,64'b1110000000000000000011000000000000000000000000000000000000000000,64'b1110000000000000000001000000000000000000000000010000000000000000,64'b1110000000000000000000110000000000000000000000111100000000000000,64'b1110000000000000000000010000000000000000000000001111100000000000,64'b1110000000000000000000010000000000000000000000000011110000000000,64'b1110000000000000000000001111100000000000000000000000011000000000,64'b1110000000000000000000000001111000000000000000000000001100000000,64'b1110000000000000000000000000011111000000000000000000001110000000,64'b1111100000000000000000000000000111110000000000000000000111100000,64'b1111111110000000000000000000000001111100000000000000000111110000,64'b1110111110000000000000000000000000000000000000000000000000110000,64'b1110001111000000000000000000000000000000000000000000000000011000,64'b1110000000111000000000000000000000000000000000000000000000011000,64'b1110000001111100000000000000000000000000000000000000000000011001,64'b1110000000011110000000000000000000000000000000000000000000001111,64'b1110000000000011100000000000000000000000000000000000000000000110,64'b1110000000000001100000000000000000000000000000110000000000000000,64'b1110000000000001100000000000000000000000000000011100000000000000,64'b1110000000000000110000000000000000000000000000000011100000000010,64'b1110000000000000010000000000000000000000000000000000000000000110,64'b1110000000000000011000000000000000000000000000000000000000000110,64'b1110000000000001011000000000000000000000000000000000000000000010,64'b1110000000000000011000000000000000000000000000000000000001111110,64'b1111000000000000011100000000000000000000000000000000000001111110,64'b1111000000000000011100000000000000000000000000000000000001111110,64'b1111000000000000001100000000000000000000000000000000000011011110,64'b1111000000000000000100000000000000000000000000000000010011010000,64'b1111000000000000110000000000000000000000000000000000011111000000,64'b1111100000000110110000000000000000000000000000000000000011111111,64'b1111110000000010000000000000000000000000000000000000000011001110,64'b1110011100000001111000000000000000000000000000000000000011111000,64'b1110000111000011111100000000000000000000000000000000000011111110,64'b1111000001111000000100000000011000000000000000000000000000110010,64'b0111111100011110010000011111111100000000000000000000001100001110,64'b0111001111001111110000000011100100000000000000000000000000000000,64'b1111000011110111110000000111111110000000000000000000000000000000,64'b1111011111111100111100000001111110000000000000000000000000000000,64'b1110011111111111111011100110011111000000000000000000000011110000,64'b0111111111111111111111111100000011100000000000000000000000000000,64'b1111111111111111111111111000001111110000111000011000000000000000,64'b1111111110011111111111111011100000111100000000000000000000000000,64'b1111111100000000000011111111110011011111100000000000000000000000,64'b1111111000000000000000011111011000000111110000000000000000000000,64'b1110000000000000000000000111111111100101111100000000000000000000,64'b1110000000000000000000000011111111110011111100000000000000000000,64'b1110000000000000000000000000111111101101111100000000000000000000,64'b1110000000000000000000000000001111111011111000001000000000000000,64'b1110000000000000000000000000000001111111111000011110000000000000,64'b1110000000000000000000000000000000011111111011010100000000000000,64'b1110000000000000000000000000000000000000000000011100000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000};
assign input_o[67] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000111110000000000000000000000000000000000000000000000000,64'b0000000001111110000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000111100000000000000000000000000000000000000000000000000,64'b0000000001111111100000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000011,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000001110000000000000000000000000000010,64'b0000000000000000000000000000000111110000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000010000000000000000000000000000,64'b0000000000000000000000000000000000011100000000000000000000000000,64'b0000000000000000000000000000000000010000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000001100000000000000000000000000000000,64'b0000000000000000000000000000000000010000000000000000001111111111,64'b0000000000000000000000000000000000010000000000000000000000111100,64'b0000000000000000000000000000000000010000000000000000000001111111,64'b0000000000000000000000000000000000000000001111111100000011111111,64'b0000000000000000000000000000000000000000111111111000000011111111,64'b0000000000000000000000000001111111000000011111111111111000000000,64'b0000000000000000000000000000000000001111111111111111111000000000,64'b0000000000000000000000000000000001001111111111111111110000000000,64'b0000000000000000000000000011111111111111100000000000000000000000,64'b1111001110000000001111000000111111110000000000000000000000001111,64'b0000111111111111111111000000000000000000000000000111111111111110,64'b1111111111111111100000000000000000000000000000000111111111100000,64'b1111111111000000000000100000000000000011111100000000000000000000,64'b1100000000000000000000100000001111111111111110000000000000000000,64'b0000000000000000000000000000001111000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000111111100000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000010000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[68] = {64'b0000000100000000000000000000000000000000000000000000000000011100,64'b0000111100000000000000000000000000000000000000000000001101111111,64'b0000000000000000000000000000000000000000000000000000000111110000,64'b0000000000000000000000000000000000000000000000000000000111000000,64'b0000000000000000000000000000000000000000000000000000001111000000,64'b0000000000000000000000000000000000000000000000000000001111000000,64'b0000000000000000000000000000000000000000000000000000001111000000,64'b0000000000000000000000000000000000000000000000000000001111100000,64'b0000000000000000000000000000000000000000000000000000001111100000,64'b0000000000000000000000000000000000000000000000000000000111100000,64'b0000000000000000000000000000000000000000000000000000000111100000,64'b0000001000000000000000000000000000000000000000000000011111111100,64'b0000001000000000000000000000000000000000000000000000011111111100,64'b0000001000000000000000000000000000000000000000000000001110111100,64'b0000001001100000000000000000000000000000000000000000001111111000,64'b0000001001100000000001000000000000000000000000000000000011111110,64'b0000001000100000000001000000000000011111111111110000000001110000,64'b0000001000100000000000000000000001111111111111111000000000000000,64'b0000001000100000000000000000000000000000111100000000000000111111,64'b0000001100100000000000000000000000000000000000000000000001111111,64'b0000001100100000000000000111110000000000000000000000000011111111,64'b0000001100100000000001001111111100000000000111100000111111111111,64'b0000000100110000000001000000000000000000001111111111111000011111,64'b0000000100010000000000000000000000000000000000001111111001111111,64'b0000000110010000000000000111000000000000001100000000000111111100,64'b0000000010010000000000000000000000000000011111111111111111110000,64'b0000000110010000000000000000000000000000111111111111111111000000,64'b0000000110000000000000000000000000000000000001111111111000000000,64'b0000000010010000000000000000000000000000000000111100000000000000,64'b0000000000010000011000000000001110000000000000000000000000000000,64'b0000000001100000000000000001111100000000000000000000000000000000,64'b0000000000010000000000000011110000000000000011100000000000000000,64'b1000000000000001111110000000011111000000000000000000000000000000,64'b0000000000000011111111000000011000000000000000000000000000000000,64'b0000000000000000000011000000100000000000000000000000000000000000,64'b0000000000000000000000111100000000000000000000000000000000000000,64'b0000000000000000000000111100000011111000000000000000000000000000,64'b0000111000000000000000000000001111111000000000000000000000000000,64'b1111111100000000000000000000011111111100000000000000000000000000,64'b0001011100000000000010000000000000001100000000000000000000000000,64'b0011001100000000011111111100001111100000000000000000000000000000,64'b0001001000000001111111111111000111110000000000000000000000000000,64'b0001101000111111111111111111110011111000000000000000000000000000,64'b0001100000000000000111111111110000000000000000000000000000000000,64'b0001100000011111111111111111110000000000000000000000000000000000,64'b1001100000000001111111111111100000000000000000000000000000000000,64'b1001000000000000000000000111100000000000000000000000000000000000,64'b0011100000000000000000001111000000000100000000000000000000000000,64'b0000001000011111000000000000000000000000000000000000000000000111,64'b0011101111111111000000000000000000000000000000000000000000111111,64'b1111111111111111100000000000000000000000000000000000000111111111,64'b1111111111111111000000000000000000000000000000000000001111111111,64'b0000111111111111111100000000000000000000000000000000001000001111,64'b0000011111111111111100000000000000000000000000000000001111111111,64'b0000001111111110000000000000000000000000000000000000001111111111,64'b0000000000000000000000000000000000000000000000000000000001111111,64'b0000000000000000000000000000000000000000000000000000000000001111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[69] = {64'b0000000000000110000000000000000000111111100000000000000000000000,64'b0000011111000010000001111111001000111111111111100000000000000011,64'b1111111100000010000000011100110111111111111110000000000000001111,64'b1111111101000011111111110000000000001111000000010000000000111111,64'b0001101011000111111111111110000000000000001111000000111110000000,64'b0000000101100011111111111000011111110000000000000011110000000000,64'b0000001111000111111111111001111111100000000000000000000000000000,64'b0100011111000000011111111111111110000110000100000000000000000000,64'b1011111000000000000000011111110000010000000000000000000000000000,64'b1100000000000111111111000000000000001111100000000000000000000000,64'b1100001111110001110001111000011100011110000000000000000000000000,64'b0000000000000000100000011000100000000000000000000000000000000000,64'b0000001000000110100000111000100000000000000000000000000000000000,64'b0000001000000110111000000000000000000000000000000000000000000000,64'b0000000000000010011000000111100000000000000000000000000000000000,64'b0000000000000111111001100011000000000000000000000000001111111111,64'b1111111111000000000000000000000000000000000000000000000000000000,64'b0001000000000000000000000000000000000000000000000000000000000000,64'b0000000000011110011100000000111000000000000000000000000000000000,64'b1111111111111111111000000000111100000000000000000000000000000000,64'b1100000001111110001000000000000000000000000000000000000000000000,64'b1111111111111111111100000000000000000000000000000000000000000000,64'b1111100000011111111000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1110001000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000011110000000000000000000000000000,64'b0000000000000000000000000000111111111110000000000000000000000000,64'b0000000000000000000000000001111111100000000000000000000000000000,64'b0000000000000000000000000000111011000000000000000000000000000000,64'b0000000000000000001000000011100011100000000000000000000000000000,64'b0000000000000000000000001100000001110000000000000000000000000000,64'b0000000000000000000100011100000011100000000000011000000000000000,64'b0000000000000000000000001111000011100000000000000000000000000000,64'b0000000000000000000000000111111001100000000000000000000000000000,64'b0000000000000000000000000111111111000000000000000000000000000000,64'b0000000000000000000000000001111111110000000000000000000000000000,64'b0000000000000000000000000000000111100000000000000000000000000000,64'b0000000000000000000000000011110000000000000000000000000000000000,64'b0000000000000000000000000001111111100000000000000000000000000000,64'b0000000000000000000000000000111111110000000000000000000000000000,64'b0000000000000000000000000000000111000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000110000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000001111111100000000000000000000000000,64'b0000000000000000000000000000011000000000000000000000000000000000,64'b0000000000000000000000000000001111111110000000000000000000000000,64'b0000000000000000000000000000000111110000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[70] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000010000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000111100000000000000000000000000000000,64'b1110000000000000000000000011111100000000000000000000000000000000,64'b1010000000000000000000000011011100000000000000000000000000000000,64'b1100000000000000000000000001111000000000000000000000000000000000,64'b1100000000000000000000000111111000000000000000000000000000000000,64'b1100000000000000000000000000001000000000000000000000000000000000,64'b1100000000000000000000000111111000000000000000000000000000000000,64'b1000000000000000000000000011110000000000000000000000000000000000,64'b1100000000000000000111110000000001111100000000000000000000000000,64'b0000000000000000000011111000000000011111110000000000000000000000,64'b0000000000000000000100000000000000000011111000000000000000000000,64'b0000000000000000000000000000000000000000011000000000000000000000,64'b0000000000000000010000000000000000000000011110000000000000000000,64'b0001111000000000111110000000000000000010000111100000000000000000,64'b0001111100000000111110000000000000000000000011110000000000000000,64'b0010001111000001111100000000000000000001111111010000000000000000,64'b0001111000000101111110000000000000000000111111100000000000000000,64'b0011111000000000011000000000000000000000000000000000000000000000,64'b0010011101100000111000000000000000000000111000000000000000000000,64'b0000111111100000111000000000000000000000011000000000000000000000,64'b0000000000000000011000000000000000000000011000000000000000000000,64'b0111111111111111110000000000000000000000011000000000000000000000,64'b0001111111101111100110000000000000000001111111000000000000000000,64'b0000011111100000000000000000000000000000011000000000000000000000,64'b0000000000000000001111111000000000000000011000000000000000000000,64'b0000000100000000000001000001111100000000011000000000000000000000,64'b0000000000000000000000100011111110000000011000000000000000000000,64'b0000000000000000000000111111111000000000011000000000000000000000,64'b0000000000000000000000000111111110000000111000000000000000000000,64'b0000000000000000000000000000000000000000111000000000000000000001,64'b0000000000000000000000000000000000000000111000000000000000000111,64'b0000000000000000000100000000000000000000111000000000000001111100,64'b0000000000000000000000000010000000000000111000000000000000000000,64'b0000000000000000000000000000000000000000111000000001111110000000,64'b0000000000000000000011111110000000000000011000011111111100000010,64'b0000000000000000000000111110000000000000011000111100011011001101,64'b0000000000000000000000000010000000000000011000001111111111111100,64'b0000000000000000000000000000000000000000011000000100000000000000,64'b0000000000000000000000100000000000000000011000000011110000000000,64'b0000000000000000000000000000000000000000010010000001111000000000,64'b0000000000000000000000000000000000000000110111000000000000000000,64'b0000000000000000000000000000000000111001000011100000000000000000,64'b0000000000000000000000011101111001111100000011000000000000000000,64'b1110000000000000000000011100000001111100001100000000000000000000,64'b1000001100000000000000111100000000111000001110000000000000000000,64'b0011111110000000000000110000000000111111111100000000000000000000,64'b1111000000000000000000110000000000000100000000000000000000000000,64'b1100000000000000000001110000000000000011111111001110000000000000,64'b0000000000000000000001110000000010011111100110000000000110000000,64'b0000000000000000000011100000001111111111111110010111111000000000,64'b0000000000000000000010000011111100111111111111100010000000000000,64'b0000000000000000000000011111111011110100000000000000000000000000,64'b0000000000000000000000000110011111110000111111110000000000000000,64'b0000000000000000000000000111111000000000100000110000000000000000};
assign input_o[71] = {64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b1100000001100000000000000000001100000000000000000000000000000000,64'b1100000000001100000000000000001110000000000000000000000000000000,64'b1100000000001000000000000000000000000000000000000000000000000000,64'b1100000000001110000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000110000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1110000011110000000000000000000000000000000000000000000000000000,64'b1100001111110000000000000000000000000000001100000000000000000000,64'b1100011111111000000000000000000000000000001000000000000000000000,64'b1100000111110000000001100000000000000000001000000000000000000000,64'b1100011111111110000000011000010000000000000000000000000000000000,64'b1100111100011010000000001100100000000000000000000000000000000000,64'b1100001000000010000000001100110000111100000000000000000000000000,64'b1100011000001110000000000010000000011000000000000000000000000000,64'b1100011000111110000000000011100000011100000000000000000000000000,64'b1100001111111110000000000000100000011000000000000000000000000000,64'b1100000111111000010000000000000000000000000000000000000000000000,64'b1100000001110000000000000000001000000000000000000000000000000000,64'b1100000001000011100000000000000110000000000000000000000000000000,64'b1100000000000000000000000000000011000000000000000000000000000000,64'b1100000000000000001000000000000001000000000000000000000000000000,64'b1100000000000000001000000000000001100000000000000000000000000000,64'b1100000000000000111110000000000000110000000000000000000000000000,64'b1100000001000000000000000000000000010000000000000000000000000000,64'b1100000010000000000000000000000000011000000000000000000000000000,64'b1100110000000000000000000000000000011000000000000000000000000000,64'b1100000000000000000000000000000000001000000000000000000000000000,64'b1101110000000000000000000000000000001000000000000000000000000000,64'b1100000000000000000010000000000000001000000000000000000000000000,64'b1100000000000000000011000000000000000011100000000000000000000000,64'b1100000000000000001010000000000000000011111000000000000000000000,64'b1100000000000000000000000000000000000000111000000000000000000000,64'b1100000000000000000000000000000000000000101110000000000000000000,64'b1100000000000000000000000000000000000000001011000000000000000000,64'b1111110000000000000000000000000000000000000111100000000000000000,64'b1100011000000000000000000011100000000000000101101000000000000000,64'b1100000110000000000000000000100000000000000011100000000000000000,64'b1100000010000000000000000000011110000000000001011000001100000000,64'b1100000000000000000000000000000010110000000000000000001100000000,64'b1100000000111100000000000000001100111100000001000000001100000000,64'b1100000000011100000000000000000001010111000000000000000000000000,64'b1110000000011100000000000000000000010001111000000000001000000000,64'b1110000000011100000000000000001000110000011111000000101000000000,64'b1110000000001011000000000001011000000000000011000011101000000000,64'b1110000000000011111111110001011000000000000000001111101000000000,64'b1110000000000000011001110001010100000000000000011111101100000000,64'b1110000000000000000000000001011000000000000000000111111000000000,64'b1110000000000000000000000010010000000000000000011111110000000000,64'b1110000000000000000000001111000000000000000000011001110000000000,64'b1110000000000000000000000011010110000000000000011100100000000000,64'b1110000000000000000000000000110010000000000000011110000000000000,64'b1110000000000000000011110000111111000000000000010111100000000000,64'b1100000000000000001000000011111111000000000000011111010000000000,64'b1110011110000000001001111100011111000000000000011111100000000000,64'b1110110000000000001000111110101111000000000000011111110000000000,64'b1111111110000000001111111110011110000000000000000000000000000000,64'b1111111111111111000011011000110010000000000000000000000000000000,64'b1100111111110110001011111000110000000000000000000000000001100000,64'b1100000000000011001101111011000000000000000000000000000011000000,64'b1100000000000011111110110010000000000000000000000000000011000000,64'b1111100000011101111101110010000000000000000000000000000001100000,64'b1100000000001001111111111111100000000000000000000000000000000000};
assign input_o[72] = {64'b0010000000000000000000000000000000000000000100000000000000000000,64'b0001110000000000000000000000000000000000000000011111110000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0001111111111100000000000000000000000000000000000000000000000000,64'b0011111111111000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000001000000000000000000000000000000000,64'b0000000000000000000000000000111111000000000000000000000000000000,64'b0000000000000000000000000000011000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000001000000000101111100000000000000000,64'b0000111111000000000000000000000000000000101000000000000000000000,64'b0011111110000000000000000000000000000011101111100000000000000000,64'b0000111000111100000000000000000000000001111111110000000000000000,64'b1111111111111000000000000000000000000111111100000000000000011111,64'b0111111111000000000000000000001000000000000000000000000000111000,64'b0000000000000000000110000011101000000000000000000000000000000000,64'b0000000000000000000000000000001000000000000000000000000000000000,64'b0000000000000000000000000000010000000000000000000000000000000000,64'b0000000000000000000000000011111110000000000000000000000000000000,64'b0000000000000000000000000011111111100000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000111110000000000000000000000000011100000000000000000000000,64'b0000000000000000000000000111000000000000000000000000000000000000,64'b0000000000000000000000001111110000000000000000000000000000000000,64'b0000000000000000000000011111110000000000000000000000000000000000,64'b0000000000000000000000000011110000000000000000000000000000000000,64'b0000000000000000000000000001110000000000000000000000000000000000,64'b0000000000000000000000000001110000000000000100000000000000000000,64'b0000000000000000000000000011111000000000000000000000000000000000,64'b0000000000000000000000000110000000000000111111110000000000000000,64'b0000000000000000000000000000000000001111111111111111000000000000,64'b0000000000000000000000000011111111111111100110000000100000000000,64'b0000000000000000000000000011111111111100000111111111110000000000,64'b0000000000000000000000000011111111111101111111111111100000000000,64'b0000000000000000000000001111111111111111111111111100000000000000,64'b0000000000000000000000011111111111110000000000000000000000000011,64'b0000000000000000000000000000000011100000000000000000000000000000,64'b0000000000000000000000000000011000000000000000000000000000000000,64'b0000000000000000000000000000011100000001000000000000000000000000,64'b0000000000000000000000000000111100000001000000000000000000000000,64'b0000000000000000000000000000111100001001000000000000000000000000,64'b0000000000000000000000000000110100001001000000000000000000000000,64'b0000000000000000000000000000110010001001000000000000000000000000,64'b0000000000000000000000000000011101001001000000000000000000000000,64'b0000000000000000000000000000001001001101100000000000000000000000,64'b0000000000000000000000000000000001001011100000000000000000000000,64'b0000000000001111100000000000010000000001100000000000000000000000,64'b1000000000000111000000000000000000000001000000000000000000000000,64'b0011100000000000000000000000000011001110000000000000000000000000,64'b0000000000000000000000000000000000000000111111111111000000000000,64'b0000000000111111111111111111111000000000000001111111100011000000,64'b1000000000000000000000011111110111111100000000000000011111111111,64'b0000000000000011111111111111111111100000000000000101000000000000,64'b0000000000000000000000000000000000000111111100011111111111111111,64'b0000000000000000000000000000000000110000000000000000011111111111,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000000000000000000000000,64'b0011000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000};
assign input_o[73] = {64'b0000000000000000000000000010000000000000000000000000000000000000,64'b0000000000000000000000000010011111000000000000000000000000000000,64'b0000000000000000000000001000000000001111110000000000000000000000,64'b0000000000000000000001111000000111100001111000000000000000000000,64'b0000011100000000000000000000000000000000000000000000000000000000,64'b1111111100000000000000000000000000000000110000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000111111000000000000000000000000000000000000,64'b0000000000000000000000101111000000000000000000000000000000000000,64'b0000000000000000000000011111000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000001111100001111000000000000000000000000000,64'b1110000000000000000000000011100000000000111000000000000000000000,64'b0100000000000000000000000011000000000011111111000000000000000000,64'b0000000000000000000000000010010001111111111111100000000000000000,64'b1111100000000000000000000010010000000101100111100000000000000000,64'b0111100000000000000000101110100000000001111111100000000000000000,64'b0000000000000000000000101000100000000000011111000000000000000000,64'b0000000000000000010000001000010000000100011111000000000000000000,64'b0000000000000000010000000000000000000000011110000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000010000000000000000000000,64'b0000000000000000000000000000000000000000010000000000000000000000,64'b0000000000000000000000000000000000000000001100000000000000000000,64'b0000000000000000000000000000000000000000001100000000000000000000,64'b0000000000000000000000000000000000000000001100000000000000000000,64'b0000000000000001000000000000000000000000000100000000000000000000,64'b0000000000000011000000000000000000000000000011110000000000000000,64'b0000000000000011000000110000000000000000000111111000000000000000,64'b0000000110000011100000100000000000000000001111111000000000000000,64'b0000000000000011100001000000000000000000001111110000000000000000,64'b0000000000000011110001000000000000000000011111110000000000000000,64'b0000000001000011100000000000000000000000011000000000000000000000,64'b0000000000000011000000000000000000000010011000000000000000000000,64'b0000000001110011000000000000000000000010011000000000000000000000,64'b1110000000000110010111111000000000000000011000000000000000000000,64'b1111111100000110011111111100000000000000011000000000000000000000,64'b1100111000000011111111111111011100000001111110000000000000000000,64'b0111100000011000000000111111011000000000001110000000000000000000,64'b0000000000000000000001111110011100100000001110000000000000000000,64'b0000000000000000001111110001100001111000001110000000000000000000,64'b0000000000000000000000000011100011111001111110000000000000000000,64'b0000000000000000000000100001101111111011111110000000000000000000,64'b0000000000000000000000000000000001111011111110000000000000000000,64'b0000000000000001111000000000011111110111111110000000000000000000,64'b0000000000000001111000000111111001111111111111000000000000000000,64'b0000000000000011111000001111111111000000010011000000000000000000,64'b0000000000000001110000011110001110111011110011000000000000000000,64'b0000000000000000110011111111111101111110000110000000011000000000,64'b0000000000000000000000101111110001000000000000001111111111111111,64'b0000000000000000010001001111000000000000000000000000000011110000,64'b0000000000000000000001110011100000000011100000000000000000011000,64'b0000000010000000000000011111111111111111111101111111111111100000,64'b0001111100000000000000101111001111111111111111111111111111111111,64'b0000000100000000000000000000000000111111111111111111111111111111,64'b0000000000000100000000011111001111111111111111111111111111111111,64'b0000001100000000000111111111111111111111111111111111111111111111,64'b0000000001101000000110011111111111100000000000000000000001111111,64'b0000000000111111110011111111110000000000000000000000000000000000,64'b0000000000111000011111111110000000000000000000000000000000000000,64'b0000000000010111111111110000000000000000000000000000000000000000};
assign input_o[74] = {64'b0000000000000000000000000000000000000000000000000000000100111100,64'b0111000000000000000000000000000000000000000000000000111111111111,64'b0000000000000000000000000000000000000000000000000000000111111000,64'b0000000000000000000000000000000000000000000000000000000111100000,64'b0000000000000000000000000000000000000000000000000000001111000000,64'b0000000000000000000000000000000000000000000000000000000111000000,64'b0000000000000000000000000000000000000000000000000000000111000000,64'b0000000000000000000000000000000000000000000000000000000111100000,64'b0000000000000000000000000000000000000000000000000000000111100000,64'b0000000000000000000000000000000000000001100000000000000111100000,64'b0000000000000000000000000000000000000000000000000000000111100000,64'b0000000000000000000000000000000000000000000000000000000111111000,64'b0000000000000000000000000000000000000000000000000000000011111000,64'b0000000000000000000000000000000000000000000000000000000111111100,64'b0000000000000000000000110000000000000000000000000000000111111000,64'b0000000000000000000000000000000111111111100000000000001111111111,64'b0000000000000000000000000000000000000000000000000000011111111110,64'b0000000000000000000000000000001111110000001000000000000011100000,64'b0000001000100000000001000001111111111111000000000000000000000000,64'b0000001000100000000000000111111111100000000000000000000000000000,64'b0000001100100000000001000101111111111111110000000000000111111111,64'b0000001100100000000000110111111111111111011110000000001111111111,64'b0000001100100000000001111111111111111111110111000000011001111111,64'b0000001100100000000011111101111000000111111111000000010011111111,64'b0000001100100000001011111100000000000011111100000000000111111111,64'b0000000110110000001001111100000000000000011110011111111111111111,64'b0000000110110000000111111100000000000000001111111111111111111000,64'b0000000110110000000111111100000000000000000111111111111111100000,64'b1000000111010000000001111100000000000000110000111111111111000000,64'b1000000111011000000001111100000011111111111100011111111100000000,64'b1000000111111000000001011100000000011111111100000000000000000000,64'b1000000111111000000000011100011111111111111100000000000000000000,64'b0000000010110000000000010000011111111111111100000000000000000000,64'b0000000001100000000000000000110000011111111100000000000000000000,64'b0000000011110000000011010000111110011111011000000000000000000000,64'b0000000000000000000000110000111110000010111000000000000000000000,64'b1000000000000000000000011111111110000010110000000000000000000000,64'b1100000000000000000000011111011110000110110000000000000000000000,64'b1100000000000001111111100000111111000110110000000000000000000000,64'b1000000000000000011111111111111000000011010000000000000000000000,64'b1100000011100110001111100111000000000011011000000000000000000000,64'b1000111100011111011111000110000000000011011000000000000000000000,64'b0111111000011101111110000000000000000001011000000000000000000000,64'b0011011000011111100111000000000000011111111100000000000000000000,64'b0011011000011101000111111110000000000011011100000000000000000000,64'b0011001111111111111111111111000000111111111100000000000000000000,64'b0011101111111111111111110111111110111111111100000000000000000000,64'b0011100111110111000111111111111110000011110000000000000000000000,64'b0001101111111111111111111111010110000000000000000000000000000000,64'b1001100011111111111111011111111100000000000000000000000000000000,64'b0001100000000000000000000111100000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000000000000000000000000,64'b0111100001111111111100000000000000000000000000000000000000000000,64'b1111000011111111111111111000000000000000000000000000000000000000,64'b1111000001111111111000000000000000000000000000000000000011111111,64'b0111110000011111111111111110000000000000000000000000000111111111,64'b0011111111111111111111111000000000000000000000000000011111111111,64'b0001111111111111111111000000000000000000000000000000011000001011,64'b0000111111111111110000000000000000000000000000000000001111111111,64'b0000001111100000000000000000000000000000000000000000001111111111,64'b0000000000000000000000000000000000000000000000000000000000000011,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[75] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000111100000000000000000,64'b0000000000000000000000000000000000000000111111110000000000000000,64'b0000000000000000000000000000000000000000111111110000000000000000,64'b0000000000000000000000000000000000000000111111110000000000000000,64'b0000000000000000000000000000000000000000000111100000000000000000,64'b0000000000000000000000000000000000000000010001111100000000000000,64'b0000000000000000000000000000000000000000010100111100000000000000,64'b0000000000000000000000000000000000000000111000101110000000000000,64'b0000000000000000000000000000000000001110000111101110000000000000,64'b0000000000000000000000000000000000111110111111111111100000000000,64'b0000000000000000000000000000000001111111111111111110000000001100,64'b0000000000000000000000000000000011111111100111111001000100111100,64'b0000000000000000000000000000000111011101111111111111111111111100,64'b0000000000000000000000000000000110111111111111111111111111111100,64'b0000000000000000000000000000000001111111100111111111111111111100,64'b0000000000000000000000000000000000000110001111111100111111011111,64'b0000000000000000000000000000000001111011111110111111111001111111,64'b0000000000000000000000000000000000000111111011111111111000000111,64'b0000000000000000000000000000000001100110000011101111111111001111,64'b0000000000000000000000000000000000000000111111100000000011000000,64'b0000000000000000000000000000000000000000011111111111111100000111,64'b0000000000000000000000000000000000000000011111000000000000000000,64'b0000000000000000000000000000000000000000011111001011111000000011,64'b0000000000000000000000000000111110000000111010000000000000000111,64'b0000000000000000000000000001111111111111111000000000000011111111,64'b0000000000000000000000000001111011111111100000000000000011111110,64'b0000000000000000000000000000011110100110001111000000000011111110,64'b0000000000000000000000000001110000111111111010000000000111111100,64'b0000000000000000000000000111110000011111111110100001111111110000,64'b0000000000000000000000000110110000000010111100100111111000000000,64'b0000000000000000000000000100000000000010011111111111100000000000,64'b0000000000000000000001000001100000000000011111111110000000000000,64'b0000000000000000000001000000000000000000101100000000000000000000,64'b0000000000000000110001110100000000000000001100000000000000000000,64'b0000000000000000011111111100000000000000000010000000000000000000,64'b0000000000000000000001111100000000000000000000000000000000000000,64'b0000000000000000000001111100100000000000000000000000000000000000,64'b0000000000000000000100111000100000000000000000000000000000000000,64'b0000000000000000000001000011011000000000001100000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000001111000000000000000000000000000000000000000000,64'b0000000000000000000001000000000000000000000000000000000000000000,64'b0000000000000011111111000000000000000000000000000000000000000000,64'b0000000000000000110000000000000000000000000000000000000000000000,64'b0000000000000011111111111000000111100000000000000000000000000000,64'b0000000000000000000000000000011001111100000000000000000000000000,64'b0000000000000000000000000000001111111000000000000000000000000000,64'b0000000000000000000000000000000011111100000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[76] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0001000000000000000000000000000000000000000000000000000000000000,64'b0001110000000000000000000000000000000000000000000000000000000000,64'b0011110000000000000000000000000000000000000000000000000000000000,64'b0000000000011000000000000000000000000000000000000000100000000000,64'b0000000000000111000000000000000000000000000000000000100000000000,64'b0000000000000001000000000000000000000000000000000000100000000000,64'b0010000000000001000000000000000000000000000000000000000000000000,64'b0010000000000001000000000000000000000000000000000000001000000000,64'b0000011000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000001111111000000000000000000000,64'b1110000000000000000000000000000000000111111111111111100000000000,64'b1111110000000000000000000000000000000111111111111111100000000000,64'b0000000000000000000000000000010000001000001000001111100000000000,64'b0000000000000011110000000000000000000001101000000000000000000000,64'b0000000000001101110000000000000000000000011110000000000000000000,64'b0000000000000011110000000000100000000000111110000000000000000000,64'b0000000000000111110000000010111100111111111111000000000000000000,64'b0000000000000011100000000110011100001111111111000000000000000000,64'b0000000000000000000000000010000011111110011110000000000000000000,64'b0000000000000000000000001010000001111110001100000000000000000000,64'b0000000000000000000000000000000000011110000000000000000000000000,64'b0000000000000000000000000000000000001110001000000000000000000000,64'b0000000000000000000000000000000111001110001100000000000000000000,64'b0000000000000000000000000000111110000111001100000000000000000000,64'b0000000000000000000000000000111111000011111100000000000000000000,64'b0000000000000000000000000001111111000011111000011000000000000000,64'b0000000000000000000000000001110111000000111010011111100000011110,64'b0000000000000000000000000001111111000000111011011111111001011110,64'b0000000000000000000000000001111111000000011011000011111111100000,64'b0000000000000000000000000001101110000000000011000000000011111110,64'b0000000000000000000000000001100100001000000000000000000000001100,64'b0000000000000000000000000000100100000000000000000000000000000000,64'b0000000000000000000000000000100000000000011000011000000000000000,64'b0000000000000000000000000000100001110000100001111111111000000000,64'b0000000000000000000000000000010000000000000000000000000000000000,64'b0000000000000000000000000000001000000100000001111111000000000000,64'b0000000000000000000000000000001111111111111111111111111000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000001100000000000};
assign input_o[77] = {64'b1111000000000000000000000000000000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1011110000000000000000000000000000000000000000000000000000000000,64'b0011000000000000000000000000000000000000111110000000000000000000,64'b1111000000000000000000000000000000000001111111111100000000000000,64'b1111111000000000000000000000000000000000000001111111000000000111,64'b1000000000000000000000000000000000000000000000000001111111111111,64'b0001110000000000000000000000000000000000000011100000011111111100,64'b0011111111100000000000000000000000000000000000000000000000000000,64'b1111111111100110000000000000000000000000000000000000000000000000,64'b1111111111101111100000000000000000000000000000000000000000000011,64'b1111111111111011111110000011110000000000000000000000000000000111,64'b1111001111111110000000001111100000000000000000000000000000000000,64'b1111111111101111111111110000011000000000000000000000000000000000,64'b1111001111111111111111100000000000000000000000000000000000000000,64'b1111001111111111111111111000110000000000000000000000000000000000,64'b1111110010001111111111111100011111111111111111110000000000000000,64'b1111110111111100000000111111100000000000000000000000000001110000,64'b1111100000000000000000011111111111111111111111000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000110000,64'b1111101100000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000110000000000000000000000000000000000,64'b1111100000000000000000000000111000000000000000000000000000000000,64'b1111100000000000000011111000010100000000000000000000000000010000,64'b1111100000000000000000111100000000000000000000000000000000001000,64'b1111100000000000000000111110000000000000000000000000000000001000,64'b1111100000000000000010011110000000000000000000000000000000000111,64'b1111100000000000000001110100000000000000000000000000000000000111,64'b1111100000000000000011100100000000000000000000000000000000000000,64'b1111100000000000000000000100000000000000000000000000000000000000,64'b1110111000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000111110000,64'b1011100111001110000000000000000001110100000000000000000000000000,64'b0011100010000000000000000000000000000000000000000000000000111001,64'b1111111011100010111111111111111111111111111111000000001111111111,64'b0111111110100000000011111111111100111111111111000000000111001111,64'b1111111111111111111111111111111111111111111111000000000000000000,64'b1111100011100000000111100000000111111111111111111111111000000000,64'b1111111111111111100011111100001111110000000000111111111111110000,64'b1111111111111111100001111000011111111111100000000000000000000000,64'b1111111111111111111100000000011111111111111111100000000000000011,64'b1111111111111100001111111100011111111111111110000000000000000000,64'b1111111111111110000000000011111111111111111111000000000000000000,64'b1111111111111110000000010100010000000000000000000000000000000000,64'b1111111111111111111111111111000000000000000000000000000000000000,64'b1111100001111111111111000000000000000000000000000000000000000000,64'b1111100000011111111110000000000000000000000000000000000000000000,64'b1111100011111111000000000000000000000000000000000000000000000000,64'b1111100000000110000000000000000000000000111110000000000000000000,64'b1111100000000000000000000000001111111111111111000000000000000000,64'b1111100000000000000000000000111111111111000000000000000000000000,64'b1111100000000000000000111111111111100011111110000000000000000000,64'b1111100000000000000000111110000000000000000000000000000000000000,64'b1111100000000000000011111111000001100000000000000000000000000000,64'b1111100000000000000000100000000000000000000000000000000000000000,64'b1111100000000000000001111110000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000};
assign input_o[78] = {64'b0000000000000000000000000000000000000000000010000000000010000000,64'b1000000000000000000000001110000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000001110000000001111,64'b0000000000000000000000000000000000000000000000000000000000001111,64'b0000000000000000000000000000000000000000000000000000000000001111,64'b0000000000000000000000000100001000000000001000000000000000001111,64'b0000000000000000000000000000001100000000001000000000000000000111,64'b0000000000000000000000000000000110000000001100000000000000000011,64'b0000000000000000000000000000000011100000001000000000000000000010,64'b0010000000000000000000000000000000000000001000000000000000000000,64'b0010000000000000000000000000000000000000001100000000000000000000,64'b0010000000000000000000000000000000000000001100000000000000000000,64'b0010000000000000000000000000000000000000011100000000000000100000,64'b0000000000000000000000000000000000000000001000000000000000100000,64'b0000000000000000000000000000000000000000001000000000000000100000,64'b0000000000000000000000000000000000000000001000000000000000100000,64'b0000000000000000000000000000000000000000000000000000000010100000,64'b0000000000000000000000000000000000000000000000000000000001100000,64'b0000000000000000000000000000000000000000000000000000000001100000,64'b0000000000000000000000000000000011111000000000000000000000000000,64'b0000000000000000000000000000000011111000000000000000000000000000,64'b0000000000000000000000000000000011111100000000000000000000000000,64'b0000000000000000000000000000000000010100000000000000000000000000,64'b0000000000000000000000000000100000110000000000000000001000000000,64'b0000000000000000000000000001100000000000000000000000110001100000,64'b0000000000000000000000000000000000000000000000000000000000100001,64'b0000000000000000000000000011000000000111110000000101000000000000,64'b0000000000000000000000000111000001111111110000110111000010000000,64'b0000000000000000000000000111000011111111110000100111001000000000,64'b0000000000000000000000000011000000001111101000111110000000000000,64'b0000000000000000000000000011001000111111100000111111010000000000,64'b0000000000000000000000000001000000000011111000000110010000000000,64'b0000000000000000000000000001011100000000000000000110010000001000,64'b0000000000000000000000000000001000011111110000000110010000001000,64'b0000000000000000000000000000001000011111111000000110111111110000,64'b0000000000000000000000000000011000011111100000000001111111111111,64'b0000000000000000000000000000111010010111100000000000111111111000,64'b0000000000000000000000000000111100100011000000000000000000000000,64'b0000000000000000000000000000111000111111000000000000000000000000,64'b0000000000000000000000000000111000111111000000000000000000000000,64'b0000000000000000000000000000001100000011000000000000000000000000,64'b0000000000000000000000000000001100000011000000000000000000000000,64'b0000000000000000000000000000001100000111000000000000000000000000,64'b0000000000000000000000000000001100000001000000000000000000000000,64'b0000000000000000000000000000000110000101000000000000000000000000,64'b0000000000000000000000000000000010000011000000000000000000000000,64'b0000000000000000000000000000000001111011000000000000000000000000,64'b0000000000000000000000000000000001001111000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000010000000,64'b0000000000000000000000000000000001110000000000000000001111111000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000001111100,64'b0000000000000000000000000000000000000000000000000000000000111000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[79] = {64'b0000000000000001000000000000000000000000000000000000000000000000,64'b0000000000000001000000000000000000000000000000000000000000000000,64'b0000000000000001000000000000000000000000000000000000000000000000,64'b0000100000000000000000000000000000000000000000000000000000000000,64'b0110110000000000000000000000000000000000000000000000000000000000,64'b0011110000000000000000000000000000000000000000000000000000000000,64'b1011110000000000000000000000000000000000000000000000000000000000,64'b0011110000000000000000000000000000000000000000000000000000000000,64'b0011110000000001000000000000000000000000000000000000000000000000,64'b0001110000000011000000000000000000000000000000000000000000000000,64'b0000100000000011000000000000000000000000000000000000000000000000,64'b0000000000000011000000000000000000000000000000000000000000000000,64'b1111000000000001100000000000000000000000000000000000000000000000,64'b0001111110000000000000000000000000000000000000000000000000000000,64'b1000001111111000000000000000000000000000000000000000000000000000,64'b0111100111111111111100000000000000000000000000000000000000000000,64'b0011111000111111111111111100000001110000000000000000001000000000,64'b0000000100000000110000000100000000000000000000000000001000110000,64'b0000000000001100000000111000000001100000000000000000001000000000,64'b0001100000000011000001111100000000110000000000000000001100000000,64'b0000000000000011111111111000000001000000000000000001101100000000,64'b0000100000000001111110000000001111000000000000000000011100000000,64'b0001100000000000111000000011111111000000000000000000011000000000,64'b0000000000000000000000000111111111100000000000000000000000000000,64'b0000000000000000000011111111001111100000000000000000000000000000,64'b0000000000000000000011111110011111111000000000000000000000000000,64'b0000000000000000000011111110100101111000000000000000000000000000,64'b0000000000000000111111111111110000010000000000101000000000000001,64'b0000000000000000111111111111111000000000000000000000000000000010,64'b0000000000000000000001111011111100000000000000000000000000000010,64'b0000000000000000000000011111111110000000000000000000000000000010,64'b0000000000000000000001001111111110000000000000000000000000000110,64'b0000000000000000000000000111111110000000000000100000000000000110,64'b0000000000000000000011001111111111000000000000100000000000000110,64'b0000000000000000000000000111111111110000000000100000000000000110,64'b0000000000000000000000000000111111110100000001100000000000000110,64'b0000000000000000000000000000110000001000111001100000000000000110,64'b0000000000000000000000000000100000010000001001000000000000000110,64'b0000000000000000000000000000000001000011010000100000000000000110,64'b0000000000000000000000000000011000111110011000100000000000000110,64'b0000000000000000000000000111000000111000001000100000000000000110,64'b0000000000000000000000001001100000000001000000100010000000000110,64'b0000000000000000000000001000110000000000000000000000000000000110,64'b0000000000000000000000000000010111000000000000000000000000100010,64'b0000000000000000000000000000000111111111111011001110000000000010,64'b0000000000000000000000000000000001111111111111000000000000000110,64'b0000000000000000000000000000000011011111111111101111000000000110,64'b0000000000000000000000000000000001111100010001111111110000000011,64'b0000000000000000000000000000000001111111111111111111000000000001,64'b0000000000000000000000000000000000011101111111100000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000011000000000000000000000000000000000000000000000000000,64'b0000000000011111100000000000000000000000000000000000000000000000,64'b0000000000000011110000000000000000000000000000000000000000000000,64'b0000000000111100011100000000000000000000000000000000000000000000,64'b0000000000001110000111100000000000000000000000000000000000000000,64'b0000000000000111100011110000000000000000000000000000000000000000,64'b0000000000000000110000111100000000000000000000000000000000000000,64'b0000000000000000000110001110000000000000000000000000000000000000,64'b0000000000000000000011000111100000000000000000000000000000000000,64'b0000000000000000000001110011111000000000000000000000000000000000};
assign input_o[80] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000001111110000000000000000000,64'b0000000000000000000000000000000000000001000000000000000000000000,64'b0000000000000000000000000000000000000000111111000000000000000000,64'b0000000000000000000000000011111000000000111110000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000001111111100000000000000000000000000000000,64'b0000000000000000000000000000000000111000000000000000000000000000,64'b0000000111111111111000001111111111111100000011100000000000000000,64'b0000000011111100000000000111001111111111110000000000000000000000,64'b0000000000000000000000000011111111111110000000000000000000000000,64'b0000000000000000000000001111100000000000000000000011111111110000,64'b0000000011110000000000000000001111100000000000000011111111110000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000001111111,64'b0000000000000111100000000000000000000000000000000000001111111111,64'b0000000000000000000000000000000000000000000000000000111111111000,64'b0000000000111111111100000000000000000000000000000000001111000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1111000000000000000000000000000000000000000011100000000000000000,64'b0000000000000000000000000000000000000000110111110000000000000000,64'b0000000000000000011111000000000000000000000101101111111111110000,64'b0000000000000000000011000000000000111111111111110000000000000000,64'b0000000000000000000100111000111111111111111111001111111100000111,64'b0000011111111110000000011111111111111110111111111110011111111111,64'b0000001111111110000000011111111110111100000000001100001111111111,64'b0000000000100000000000001110011110111100000000000000000000111111,64'b0000000000000000000000001111111111111100000000000000000011111111,64'b0000000011000000000000000001111111111000000100000011111111111111,64'b0000001111111100000100000000000000000000111111110000000111101111,64'b0000000000000000000100000000000000000000000000000011111111111111,64'b1110000001111111111100000000000000000000000000000000000001110000,64'b1111111111111111111000000001110000000000000000000000000001000000,64'b1111111111000000000011111111110000000000000000000000000000000000,64'b1111111101111111111111111110010000000000000000000000000000000000,64'b0000000000111111111110000000000000000000000000000000000000000000,64'b0000000000000000000000000000100000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000001111,64'b0000000000000000000000000000010000000000000000000000000000000000,64'b0000000000000000000000000111110000000000001111100000000000011111,64'b0000000000000000000000111111000000000000000000000000000000001111,64'b0000000000000001111100111000000000000000000000000000000000000000,64'b0000000000000000000000000001110000000000000000000000000000000000,64'b0000000000000000111100000000000000000000000000000000000000001111,64'b0000000000000000000100000000000000000000000000000000000000111111,64'b0000000000000000001111000000000000000000000000000000000000001111,64'b0000000000000011111100000000000000000000000000000000011111111111,64'b0000000000000000000000000000000011111111111111111111111111110111,64'b0000000000000000000000000000000001111111111111111110011111111011,64'b0000000000001100000111111111111110001111111111111111111111111111,64'b1111111111111111111111100000001100000000111111111111111100000100,64'b1111111111111111100011111111111111110000000000000000000000000000,64'b1111111111000000000011111111111111111111000000000000000000000000,64'b1111111111111111110000000000010110000000000000000000000011111110};
assign input_o[81] = {64'b0000000000000000000000000000000000000000001000111100000000000000,64'b0000000000000000000000000000000000000000001000001110000011111111,64'b0000000000000000000000000000000000000000001000001000000011111111,64'b0000000000000000000000000000000000000000001000001000000000011111,64'b0000000000000000000000000000000000000000001000000000000100111010,64'b0000000000000000000000000000000000000000001000000000101100111111,64'b0000000000000000000000000000000000000000001011100000100000111110,64'b0000000000000000000000000000000000000000011110001000000000111110,64'b0000000000000000000000000000000000000000001110001000000000011010,64'b0000000000000000000000000000000000000000001110001000000000011110,64'b0000000000000000000000000000000000000000001110000000000000000100,64'b0000000000000000000000000000000000000000001110001000000000000000,64'b0000000000000000000000000000000000000000000000001000100000000000,64'b0000000000000000000000000000000000000001100000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000011111000000000001000000000,64'b0000000000000000000000000000000000000000000110000000001100000000,64'b0000000000000000000000000000000000000000001110000000001100000000,64'b0000000000000000000000000000000000000000001110000000001100000000,64'b0000000000000000000000000000001100000000001000001000000110001000,64'b0000000000000000000000000000111111100000000000001100000110000000,64'b0000000000000000000000000000111111110000000000001000000100000000,64'b0000000000000000000000000000110001111000000000000011111000000000,64'b0000000000000000000000000000110011111100000000000011111000000000,64'b0000000000000000000000000000110011111100000001000000000000000000,64'b0000000000000000000000000000110010011100000000000000000000000001,64'b0000000000000000000000000000110000011100000000000010111100000011,64'b0000000000000000000000000000110000011110001111000000000000000000,64'b0000000000000000000000000000110000001110011111001100000000000000,64'b0000000000000000000000000000110000001100111111001101111000000111,64'b0000000000000000000000000000110000100111101001001111111111111111,64'b0000000000000000000000000000110001100011100110001111111111111111,64'b0000000000000000000000000000110001110011001111111111111111110110,64'b0000000000000000000000000001110001111011000111111101111111111111,64'b0000000000000000000000000001110001111111100000001100011111111111,64'b0000000000000000000000000001100001111110000000001100011111111111,64'b0000000000000000000000000001000000111110000000000011111111111111,64'b0000000000000000000000000001000000001111000000000011111111111111,64'b0000000000000000000000000001000000001110000000000000111111111110,64'b0000000000000000000000000001000010001110000000000000000000000000,64'b0000000000000000000000000000000010000110000000000000000000000000,64'b0000000000000000000000000000000110001111000000000000000000000000,64'b0000000000000000000000000000001111111111000000000000000000000000,64'b0000000000000000000000000000000011100011100000000000000000000000,64'b0000000000000000000000000000000011111001111100000000000000000000,64'b0000000000000000000000000000000000111100111110000000000000000000,64'b0000000000000000000000000000000000111111100111000000000000000000,64'b0000000000000000000000000000000000000111111001000000000000000000,64'b0000000000000000000000000000000000000001111110000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[82] = {64'b0100000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000011110000000000000000000000000111111110000000,64'b0000000000000000011111000000000000000001111110000001111111111111,64'b0000000000000000000111100000000000000011111100011111110000000000,64'b0011110000000000000000000000000000000001111110000111111111111111,64'b0000000000000000000000000000000000000000000000001111100000011111,64'b0001000000000000000000000000000000000000000000000011110000111111,64'b0000000000000000000000000000000000000000000000000000000000111111,64'b1100000000000000000000000000000000000000000000000000000000011111,64'b1110000000000000000000000000000001111111110000000000000000000011,64'b1110000000000000000000000000000010000000000000000000000000000000,64'b0100000000000000000000000011100000111111000000000000000000000000,64'b0000000000000000000001100000000001111110000000000000000000000000,64'b1111100000001111000000001111111101111000000000000000000000000000,64'b0000000000000000000000000011111010010000000000000000000000000000,64'b0000000000000000000000000000000011111110000000000000000000000000,64'b1000000000011111000000000000000011111110000000000000000000000000,64'b1110111110111111111100001110000010111100000000000000000000000000,64'b1111111111111111111100100011111000111100000000000000000000000000,64'b1111000011100000000000100000001100000000000000000000000000000000,64'b0000000000000000000000111000000000000110000000000000000000000000,64'b0000000000000000000011110000000001111111100000000000000000000000,64'b0000000000000000000111111111000000111111100000000000000000000000,64'b0000000000000000000111111111100000000111100000000000000000000000,64'b0000000000000000001111111101000000001011100000000000000000111111,64'b0000000000000000001111011110000000001011100000000000001000111111,64'b0000000000000000001111100000000000001111100000000000000111000000,64'b0000000000000000001111010000000000001111100000000000011111111111,64'b0000000000000000001111100000000000001111100000000000000111011111,64'b0000000000000000000011110000000000000111100000000000000011111111,64'b0000000000001000010011101000000000001110100001111111111111111111,64'b0000000000000100100011100000000000001000100000000000000000000000,64'b0000000001111100000011100000000000111000101000000000000000000011,64'b0000000000000010001011100000000000111110111000000000000000000000,64'b0000000000111111111011100000000000011111100000000000000000000000,64'b0000000000000000111111100000000000010001110000000000000000000000,64'b0000000000000001111000110110110110111111000000000000000000000000,64'b0000000000000000000001111011110110100001100000000000000000000000,64'b0000000000000000000001111111111111100000000000000000000000000000,64'b0000000000000000000001111111111111100000000000000000000000000000,64'b0000000000000000111111111111001111100000000000000000000000000000,64'b0000000000001001111111111111001111100111110000000000011111111111,64'b0000000000000000111111111111001100000000000000000011111111100000,64'b0000000000000000011111111111101000000000000000000000111111111111,64'b0000000000000000011100001111100001110000000000000000000000011111,64'b0000000000000000011000101111100010100000000000000000000000000000,64'b0000000000000000011000110111100111110000000000000000000000000000,64'b0000000000000000000000101101110000100000000000000000000000000000,64'b0000000000000000000000001111100000000000000000000000000000000000,64'b0000000000000000000000000111100000000000000000000000000000000000,64'b0000000000000000000000001111100000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[83] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000011111000000000000000000000000000111111,64'b0000000000000000000000000000000000000000000000000000001111100000,64'b0000000000000000000000000000000000000000000000000000000100000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000001111000000000000000000,64'b1111111110000000000000000000000000000000011111000000000000000000,64'b0000000001000000000000000000000000000000011000000000010000000000,64'b0000000000001100000000000000000000000000000111110000010000000000,64'b0000000000000000000000000000000000000000000111111000000000000000,64'b0000000000000000000000000000000000000000000011110000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000111100000000000,64'b1111111111111100000000000000000000000000000000000011110000000000,64'b1111111111111111111000000000000000000000000000001111111111111000,64'b1111111111111111000000000000000000000000000000001111111111110000,64'b1111111111100000000000000000000000000000000000000000000000000000,64'b1111111111111100000000000000000000000000000000000000000000000000,64'b1111111111111000000000000000000000000000000000000011111111000000,64'b0000000000000000000000000000011100000000000000000000000000000000,64'b1111000001000000000000000000011111111000000000000000000000000000,64'b0011000001000000000000000000000000000000000000000111111111100000,64'b0011000000000000000000000000000000000000000000000000000000000000,64'b0011000000000000000000000000000011111100000000000111111111111000,64'b0010000001000000000000000000000000011000000000000111111000000000,64'b0010000001000000000000000000000000000000000000011000000000000000,64'b0000000000000000000000000000000000000000000000000011000000000000,64'b0000000001000000000000000000000000000000000000000110000000000000,64'b0000000000000100000000011111111100000011110000000000000000011111,64'b1111111110110100000000000111111111000000000000000000000000000000,64'b0011000000000100000000001111110111000000000000000000000000000000,64'b0001100000000100000000011100000010000000000000000000000000000000,64'b0001000000000100000000001111111000000000000000000000000000000000,64'b0000000000000100000000001111110000000000000000000000000000000000,64'b0000000000000100000000000110000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0001000000000000000000000000000000000000000000000000000000000000,64'b0001000000010000000000000000000000000000000000000000000000000000,64'b0001000000000000000000000000000000000000000000000000000000000000,64'b1001000000000000000000000000000000000000000000000000000000000000,64'b0001000000000000000000000000000000000000000000000000000000011111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000001101111111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1111100000001100000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1111111110000000000000000000000000000000000000000000000000000000,64'b1111111110000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[84] = {64'b0000001110100000010010000000000000000000100000000000000000000000,64'b0000111111110111111110111111111111111111000000000000000001111111,64'b1111111111111111110010011111111111100000000000000000011111111111,64'b1111111111111111111111111100000000000001100000011111111111111111,64'b0000000000000000000001110011111111111100000000000011000001100000,64'b0000000000111111111111111111111111100000000000000011111111111111,64'b0000000111111111111111111111111111110000000000000011111111100000,64'b0001111111111111111111111111101111111110000000000000000000000000,64'b0011111111111111111111111111111111111000000000000000000000001111,64'b0001111101111111111111111111111111111100111110000000000000000111,64'b1110011111111110000000000000000011100111111100000000000100100011,64'b1000000011100000010000000111111111111111000000000000000001111111,64'b0010000000011111111000001111111111111111000000000000000000000000,64'b0010000011111111100000111100001100100011100000000000101111111111,64'b0010111111111101100000111000100011111000100000000000111111111111,64'b0011111111111111100000100000011111111111111111111110110000000000,64'b1111111111111111000001111000100000000000011111111000000000000000,64'b1111111111111100000000111101111111111000001000000000011111111111,64'b1110001111110000000000111111111000000000000000000000111111111111,64'b0000000000000000000000110011111111111100000001111100001111111111,64'b1111111111111111111111110111111111111110001111111110100000111111,64'b1111111111111111111110000000000000000000100000000001111111111111,64'b1111111111111111111000000000000000000000000111111110001111110000,64'b1111111111111111000000000000000000000000001111111111111111111111,64'b1111111111111111000000010000000000000000000000000000110111111111,64'b0000000000000000000000011000000000000000000000000000110000111111,64'b0000000000000000000000010000000000000001001111111111100000000000,64'b0000000000000000000000010001100000000000001111111111111111110000,64'b0000000000000000000011110010010111001110101111001111110011111111,64'b0000000000000000000000000000000000000000001111100110001111111111,64'b0000000000000000000000000000000000000000000111111111111111110000,64'b0000000000000000000000000000100000000000000000000011111111111111,64'b0000000000000000000000000000100000000000000000000000011111111111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000001100100000000001,64'b0000000000000000000000000000000000000000000000000110100001111111,64'b0000000000000000011000000000100000000000000000000001111100011111,64'b0000000000000000000000000000100000000000100000000000111001111111,64'b0000000000000000000000000000100001000000100000000000111000001010,64'b0000000000000000000000000000000000000000100000000000111100000010,64'b0000000000000000000000000000010000000000100000000000001110000111,64'b0000000000000000000000000000000000000000000001111111100110001111,64'b0000000000000000000000000000010000000000001111111111111000000111,64'b0000000000000000000000000000000000000000000000011110011100000011,64'b1100000000000000000000000000000000000000000000000000001111110111,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b0001000000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000001111111111100000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b0000100000000000000000000000000000000000011111111111110000000000,64'b1000100000000000000000000000000000000000000111111111000000000000,64'b1111111111000000000000000000000000000000000000000000000000000000,64'b1111111111100000000000000000000000000000000000000000000000000000,64'b1111111111000000011111111111111111111111110000000000000000000000,64'b0001000000011100000000110011111100000000000001111100000000000000,64'b0001100111111111111100011111111111111100011111111100000000000000,64'b0000011111100001111111111111111111111111100000001111100000000000,64'b1111111111111111111111111111111111111111111111111111000000000000,64'b0001100111111111111111110000000000011111111111111111110000000000,64'b1111100000000000000000000000000000000000000000000000001100000000,64'b1111111000000000000000000000000000000000000000000001111111000000,64'b0000000000000000000000000000000000000000000000000000000001111111,64'b0000000000000000000000000000000000000000100011111111110000011111};
assign input_o[85] = {64'b0000000000000000000000000000000000000000000000000000001000000000,64'b0000000000000000000000001110111110000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000111000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000010000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000001111111111111111111111,64'b0000000000000000000000000000000000000000000000000000000000011110,64'b0000000000000000111000000000000000000000111111111111111111111110,64'b0000000000000001100000000000000000000011111111111111111111111111,64'b1111111111111111000000000000000000000000000000000000000000000000,64'b1111111111110000000000000000000000000000000000000011110000000111,64'b1111111111000001100000000000000000000000000000000000000000000000,64'b0001111111100000110000000000000000000000000000000011111100000000,64'b1111111111111111111100000000000000000000000000000000000000000000,64'b1111111111111100000000000000000000000000000000000000000000000000,64'b1111111110000000000000000000000000000000000011000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000111111,64'b0000000000000000000000000000000000000000000000000000000001111111,64'b0000000000000000000000000000000000000000000001110001111111111111,64'b0000000000000000000000000000000000000000001111111111111111100001,64'b0000000000000000000000000000000000000000011111111111111111000000,64'b0000000000000000000000000000011111111111111110000010011111100000,64'b0000000000000000000000000000111111111111110000111111111111000000,64'b0000000000000000000000000111000000000000000011111111111000000000,64'b0000000000000000111111111111100000000000000111111100000000000000,64'b0000000000000001111111111111111110000000000000000000000000000000,64'b0001111111111111111111100000010000000000010000000000000000000000};
assign input_o[86] = {64'b0000000000000000000000000000000000000000010100000000100000000000,64'b0000000000000000000000000000000000000000111000000000100000000000,64'b0000000000000000000000000000000000000000111000000001100000000000,64'b0000000000000000000000000000000000000000111000000001000000000000,64'b0000000000000000000000000000000000000001010000000001000000000000,64'b0000001111111110011111100000000000000101110000000000000000111111,64'b0000100000000011110000000000000000000011100000000010000000000000,64'b0000000000011111100110000000000000000011100000000100000000000000,64'b0000000000011111111111111000000000000111000000000100000000000000,64'b0000100000111111111011111111111111000101000000000100000000000000,64'b0000001110011001111110011111110110101111000000000100000000000000,64'b0000000001111000000000111100001111001010000000000000000000000000,64'b0000000000001100000000001110010001110110000000000000000000000000,64'b0000000000000110010000111100000000110100000000000000000000000000,64'b0000000000000011101111111000010010000100000000000000000000000000,64'b0000000000000001111111101111111111100100000000000000000000000000,64'b0000000000000000011100000111111111111110000000111000000000000000,64'b0000000000000000011110011011111100000011000000011000000000000000,64'b0000000000000000111000000001101101000011100000000000000000000000,64'b0000000000000000110000000001111100110111110000000000000000000000,64'b0000000000000001111000000000000000000001110000000000000000000000,64'b0000000000000011100000000000000000000001110000000000000000000000,64'b0000000000000111000000000000000000001111110000000000000000000000,64'b0000000000000111000000000000000000000110000000000000000000000000,64'b0000000000000111000000000000000000000110000000000000000000000000,64'b0000000000000011000000000000000000000011000000000000000000000000,64'b0000000000000001110000000000000000000011000000000000000000000000,64'b0000000000000001110000000000000000000011000000000000000000000000,64'b0000000000000000111100000000000000001011000000000000000000000000,64'b0000000000000000010010000000000000001011000000000000000000000000,64'b0000000000000000010000001111000000001001101000000000000000000000,64'b0000000001111111111111011111000000001001101000000000000000000000,64'b0000000001001010000000101011000000000001100000000000000000000000,64'b0000000000111111111111100110000000000000110000000000000000000000,64'b0000000000000000011111111111100000000000110000000000000000000000,64'b0000000000000000111000001111000000000000011000000000000000000000,64'b0000000000000000111100110000000000000000011000000000000000000000,64'b0000000000000000011000000000000000000000011000000000000000000000,64'b0000000000000000011100000000000000000000111000000000000000000000,64'b0000000000000000011000000000001110000101110000000000000000000000,64'b0000000000000000011100000000001111111111110000000000000000000000,64'b0000000000000000110110010000101111101001000000000000000000000000,64'b0000000000000000011111101111111111100011111000000000000000000000,64'b0000000000000000000101111111111001111001110110000000000000000000,64'b0000000000000000001110111111000000111100011011000000000000000000,64'b0000000000000000111011111111000000000011111110000000000000000000,64'b0000000000000000011101000101100000000011111111010000000000000000,64'b0000000000000000101111101011100000000000001101101000000000000000,64'b0000000000000111111101110011000001000000001000110000000000000000,64'b0000000000001111110111110010000001000000001111111000000000000000,64'b0000000000011111110111000010000000000000000011111000000000000000,64'b0000000000000111110111100111000000000000000001101100000000000000,64'b0000000001101110000110111111111110000000000000010111100000000000,64'b0000000000001010000000001111000000000000000000001111101000000000,64'b0000000000001000000000000111011100000000000000000110111100000000,64'b0000000000011000000000001111111000000000000000001011011100000000,64'b0000000000011000000000000000000000000000000000000000011000000000,64'b0000000000111000000001010000000000000000000000000000011000000000,64'b0000000000111000000011000000000000000000000000001110000000000000,64'b0000001111111000000000000000000000000000000001000110000000000000,64'b0000000110111000000000000000000000000000000001110100000000000000,64'b0000011111101000000000000000000000000000000001000100000000000000,64'b0001111111000000000000000000000000000000000111000000000000000000,64'b0000111011000000000000000000000000000000000000000000000000000000};
assign input_o[87] = {64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000011000000000,64'b1110000000000000000000000000000000000000000000000001100000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000011100000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000011111000000000000000000000000000000000000000000000,64'b1110000000001111111110000000000000000000000000000000000000000001,64'b1110000000001111111110000000000000000000000000000000000000001111,64'b1111000000001111110110000000000000000000000000000000000000000011,64'b1111000000000111100100000000000000000000000000000000000000000000,64'b1111000000100011100001001111111000000000000000000000000000000000,64'b1111000000000001111111111111111110000000000000000000000000001110,64'b1111000000000000011000000000011111100000000000000000000000000000,64'b1111000000000000110000000000111111111000000000000000000110000000,64'b1111000000001000110000000000011101111000000000000000000000001110,64'b1111000000001000110000000000001111011100000000000000001111111000,64'b1111000000100000110000000000000011101110000000000000011100000000,64'b1111000000110000110000000000010000110110000000000011100000110011,64'b1111000000110000010000000000000000001111000000010000000000111000,64'b1111000000100001110000000000100000000101110000100000000000000111,64'b1111000000100001111110000000000000000101110000000000000001111100,64'b1111000000101001100001000000000000000000110000000000000111000000,64'b1111000000100000110000000000000000000101111000000000111000000000,64'b1111000000100111110100000000000000000000110000011110000000000000,64'b1111000000000000111011000000000000000011110000111000000000000000,64'b1111000000001111011111000000000000000000011110000000000000000000,64'b1111000000000010011111111100000000000000011110000000000000000000,64'b1110000000000000000111110000000000000000011111100000000000000000,64'b1110000000000000000111100011000000000000011111000000000000000000,64'b1111000000000000001111111101000000000000000111110000000000000000,64'b1111000000000000000011111111100000000000111111100100000000000000,64'b1111000000000000000111010001111000000111111101100110000000000000,64'b1111000000000001111110110110010000000101111111111100000000000000,64'b0110000000001111100110111010001000000111011111111100000000000000,64'b1110000001111100000000001000001010111101110111111100000000000000,64'b1110000111100000000000000110111010001110010111100000000000000000,64'b1111110000000000000000000000011000110111100110000000000000000000,64'b1111000010000000000000000000000111110011111110000000000000000000,64'b1110000000000000000000000000001111110001111111100010000000000100,64'b1110000000000000000000000000000111111011111111100000000000001000,64'b1110000000000000000000000000000111101110111101110110000000000000,64'b1110000000000000000000000000000001111111011111110000001111000000,64'b1110000000000000000000000000000000111111101111110000111100000000,64'b1110000000000000000000000000000000011111110111111111111110000000,64'b1110000000000000000000000000000000011111111001111110010000000000,64'b1111000000000000000000000000001111111111111111111011001110000000,64'b1111000000000000000001100001111100000001111111111111000000000000,64'b1111000000000000000000111110000000000001111111111010000000000000,64'b1110000000000000000000000000000000000000111111110110110000000000,64'b1110000000000000000001000000000000000001001111011111111000000000,64'b1110100000000000000000000000000000000000000011111110110000000000,64'b1110011000000000000000000000001110000000000001111111101111000000,64'b1111110001111110000000000000111100000000000000011111111111111110,64'b1110011110000000100000000000000000000000000000001111110111111111,64'b1110000000100000000000110000000000000000000000000001111111111100,64'b1110000000000000001111110000000000000000000000000000011111110101,64'b1111000000000011111100000000000000000000000000000000000111100000,64'b0111000000011111100000000000000000000000000000000000000011100000};
assign input_o[88] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000011111100000000000111,64'b0000000000000000000000000000000000000000000000111100000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000111111111,64'b0000000000000000000000000000000000000000000000000000000011111111,64'b0000000000000111110000000000000000000000000000001110000000000111,64'b0000000000011111111000000000111100000000000000000000011000000000,64'b0000000000011111110000000000111110000000111111111111111111111111,64'b0000000000011111110000000111111111100000001111111111111111111111,64'b0000000000011011110000000111111111100000000000000000000000111111,64'b0000011111110011000000000111100011111000111100000000000000000000,64'b0000111111110011000000000111111101111000000000000000000000000000,64'b0000111100001111110000000000110100111000000000000000000000000000,64'b1000110000011111111100000000011000111000000000000000000000000000,64'b1111000000011111111110000000011000111100000000000000000000000000,64'b1111100000001111011110001111001000111110000000000000000000000000,64'b1011100000000111111110000000010011100111100000000000000000000000,64'b1110000000000011111100000000000111111111110000000000000000000000,64'b1110011110000000000000000000000000011111111000000000000000000000,64'b1111111111111000000001100000011110001111111000000000000000000000,64'b1111100000111000000011100011100000001110111000000000000000000000,64'b1111000000000011100001100011100100011101111000000000000000000000,64'b1110000000000000000111100011101111111111111000000000111000000000,64'b1100011100000000000000000001110000100111111100000001111111100000,64'b1111000000000000000000000000000100001110011111000001111111111000,64'b1110010000000111000000000000000000010011001111000011111111111110,64'b1110000000000000000000000000000000000000000111000001111101111111,64'b1110000000000000000000000000000000000000000000111110011111001111,64'b1111110000000000000000000000000000000000000000111111000111100111,64'b0001110000000000000000000000000000000000000000000011111000000000,64'b0111000000000000000000000000000000000000000000011011111111000000,64'b1111000000000000000000000000000000000000000000000111111111111101,64'b1111111100000000000000000000000000000000000111111001111111000000,64'b1111100000000000000000000000000000000000000000000000001111100000,64'b1111110000000000000000000000000000000000000000000000000111111000,64'b1110010000000000000000000000000000000000000000000000000000000000,64'b0000010000000000000000000000000000000000000000000000000000000000,64'b0000010000000000000000000000000000000000000000000000000111111000,64'b0001110000000000000000000000000000000000000000000000000011000000,64'b0111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1110110000111111111110000000000000000000000000000000000000001111,64'b1000000001111111001111110000000000000000000000000000000001111101,64'b0000011111111111111111111000000000000000000000000000000010001111,64'b1000011111111111111111000000000000000000000000000000000011111111,64'b1110000111111111110000000000000000000000000000000000000111111111,64'b0110000000000000010111110000010000000000000000000000000111111000,64'b1100010111111110000000000000111000000000000000000000000111000000,64'b1001110001111111000000000001111000000000000000000000000111000000,64'b0001110000000000000000000111111000000000000000000000000111000000,64'b0000000000010000001111111111111000000100000000000000000111100000,64'b0000000000001100011111100111111010000000000000000000000111100000,64'b0000000000001110011111100101111100000000000000000000000001110000};
assign input_o[89] = {64'b0000000000000000000010000000110000000000000000101000000000000000,64'b0000000000000000000000000001000001100000000000000000100000000000,64'b0000000000000000000000000000011111110000000000011000011111000000,64'b0000000000000000000000000000011101110000000000001000000000000000,64'b0000000000000000000000000000001111110000000000000011111100000000,64'b0000000000000000000000000000001111110000000000000000000000000000,64'b0000000000000000000000000000000100110000000000000000011111111110,64'b0000000000000000000000000000000000100000000000000000001111111110,64'b0000000000000000000000000000000001000000000000000000001111111110,64'b0000000000000000000000000000001111100000000000000000111111111100,64'b0000000000000000000000000000000000000000000000000000000000011000,64'b0000000000000000000000000000000000000000000000000000000000010000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000011111100000000000000000000000000000,64'b0000000000000000000000000000111111100000000000000000000000001110,64'b0000000000000000000000000000111111100000000000000000000000011111,64'b0000000000000000000000000000111111100000000000000000000000000000,64'b0000000000000000000000000000011101111100000000000000000000000000,64'b0000000000000000000000000111111111111111100000000000000000000000,64'b0000000000000000000000001111111101101111111000000000000000000000,64'b0000000000000000000000111111000000000001111100000000000000000000,64'b0000000000000000000001110000000001111110111100000000000000000000,64'b0000000000000000000001111000000000000000011110000000011111100000,64'b0000000000000000000011001100000000000000001110000011111111110000,64'b0000000000000000000011000110000000000000001111101111111111110000,64'b0000000000000000000110000111100000000001110011111111001111110000,64'b0000000000000000000110000100000000000000111101111000000101110000,64'b0000000000000000000110100110000000000000011111111101111111110000,64'b0000000000000000000111101100000000000011111111101110111111110000,64'b0000000000000000000111100000000000011111111011111111111111111000,64'b0000000000000000001110100010000000000011111000111111111111100000,64'b0000000000000000001110000011100000000000011100000111111000000000,64'b0000000000000000001111110011000000000111111100000000001111110000,64'b0000000000000000001110110011110000011111111100000000101111111110,64'b0000000000000000000111111111111111111111111100000000100011100000,64'b0000000000000000000011111111101100000001111000000000100000010010,64'b0000000000000000000000000001110111111011111100000000110000000000,64'b0000000000000000000000000000111110011011100000000000111110011110,64'b0000000000000000000000000000110000011011100000000000111000111110,64'b0000000000000000000000000000110000111111100000000000011000101110,64'b0000000000000000000000000000111010011111100000000000011000101110,64'b0000000000000000000000000000011010011111100000000000011000101110,64'b0000000000000000000000000000011010011111100000000000011000101110,64'b0000000000000000000000000000011000011111100000000000011000101100,64'b0000000000000000000000000000011000011111100000000000011000101100,64'b0000000000000000000000000000011000000111100000000000011000101100,64'b0000000000000000000000000000011000000111100000000000011111101100,64'b0000000000000000000000000000001000000001100000000000011000101100,64'b0000000000000000000000000000001111100110001000000000000111111010,64'b0000000000000000000000000000001101100001000000000000001111111111,64'b0000000000000000000000000000000111111111111100000000000111011110,64'b0000000000000000000000000000001111111100000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[90] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000011111100000000000000000000000011111111100000000,64'b1111111111111111111111111111111111110011110001110000000000000000,64'b1111111111111111111111111111111111111111111111111111111111000000,64'b0000000000000100000000000000000000000000000000000000000000000000,64'b1111111111111111111111111111111111111111111111111111100000000000,64'b1100000011111111000001111000000000000000000000000000000000000000,64'b0000000000111110000000111111110000000000000000000000000000000000,64'b0000000000000000000000000011110000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0001110000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1100000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000001110000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000111110000000000000000000000000000000000000,64'b0000000000000000000000111000001100000000000000000000000000000000,64'b0000000000000000000000101111100000000000000000000000000000000000,64'b0000000000000000000000001100000000000000000000000000000000000000,64'b0000000000000000000000000000000001000000000000000000000000000000,64'b0000000000000000000000000000011111000000000000000000000000000000,64'b0000000000000000000000000001111110110000111110000000000000000000,64'b0000000000000000000000000001110000000001111111000000000000000000,64'b0000000000000000000000000001100000010111111111000000000000000000,64'b0000000000000000000000000001100000000000000000000000000000000000,64'b0000000000000000000000000000100000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000111000000000000,64'b0000000000000000000000000001111111000000000000000111000000001000,64'b0000000000000000000000000011111101000000000000000111000000000000,64'b0000000000000000000000000100111111111000000000000000000000000000,64'b0000000000000000000000000001101111011111110000000000000000000000,64'b0000000000000000000000000001111111111111111000000000000000000000,64'b0000000000000000000000001001011100111111111100000000000000000000,64'b0000000000000000000000001100111000011111111111110000000000000000,64'b0000000000000000000000001100001000000111111100000000000000000000,64'b0000000000000000000000000111111111000001111111000000000000000000,64'b0000000000000000000000000110011000000000111100000000000000000000,64'b0000000000000000000000000011110000000000000000000000000000000000,64'b0000000000000000000000000000100000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000111111110000000,64'b0000000000000000000000000000000000000000000000111111111110000000};
assign input_o[91] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000110000000001110000000,64'b0000000000000000000000001110000000000000000000000100011111110000,64'b0000000000000000000000000000000000000000000100001011100000000000,64'b0000000000000000000000000000000000000000001111111011100000000000,64'b0000000000000000000000000000000000000001011111111011000000000000,64'b0000000000000000000000000000000000000001111100000111000000000000,64'b0000000000000000000000000000000000000000111100000011000000000000,64'b0000000000000000000000000000000000000000011100101101000000000000,64'b0000000000000001111111000000000000000000011111101000000000000000,64'b0000000000000111111111110000000000000000000111111000000000000000,64'b0000000000111111111011110000000000000000000000000000000000000000,64'b0000000000111111111111110000000000000000000000000000000000000000,64'b0000000000110100000001110000000000000000000000000000000000000000,64'b0000000000010010001111110000000000000000011111111000000000000000,64'b0000000000110000000111110000000000000000011110110000000000000000,64'b0000000000110000001001111000000000000000001111110000000001111000,64'b0000000000111001000011011000000000000000000011111000000000000000,64'b0000000001111000001111110000000000000000000000000000110000000000,64'b0000000001111000011100000011100000000000000000000000100000000000,64'b0000000011110000000011100011111100000000000000000000000000000000,64'b0000000011000000000001110001001111000000000000000000000000000000,64'b0000000011000000000011100001110011100000000000000000000000000000,64'b0000000011100000000000000000000001111000000000000000000000000000,64'b0000000001100000000000000000000000011000000000000000000000000000,64'b0000000000110000000000000000000000001110000000000000000000000000,64'b0000000000111000000000000000000000000011100000000000000000000000,64'b0000000000011000000000000000000000000011000000000000000000000000,64'b0000000000011000000000000000000000000000000000000000000000000000,64'b0000000000011000000000000000000000000000100000000000000000000000,64'b0000000000001100000000000000000000000000100000000000000000000000,64'b0000000000011000000000000000000000000000000000000000000000000000,64'b0000000000001100000000000000000000000000011111111000000000000000,64'b0000000000001100000000000000000000000000011111111001000000000000,64'b0000000000001100000100000000000000000000000111111001000000000000,64'b0000000000001100000100011000000000000000000011111111000000011000,64'b0001000000000110000010000110000000000000000011111100000000001000,64'b0110000000000110101000110001100010000000000000011000000000000000,64'b0100000000000010000011111000000000000000000000000000000000000000,64'b0000000000000000111001011110111110000000000000000000000000000000,64'b0000000000000000110011111111111111100000000000000000000000001000,64'b0000000000000000111111101111111110000000000000000000000000001000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000010000000000000000000000000000000000000,64'b0000000000000000000000000010000000000000000000000000000000000000,64'b0000000000000000000000000000011100000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000001110000000000,64'b0000000000000000000000000000000000000000000001100011110000000000,64'b0000000000000000000000000000000000000000000000011100110000000000,64'b0000000000000000000000000000000000000000000111111001110000000000,64'b0000000000000000000000000000000000000000000000001100000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[92] = {64'b0100000000000000000000000000000000000000000001000000000000000000,64'b0111000000000000000000000000000000000000001100100000000000000000,64'b1011100000000000000000000000000000000000000000010000000011000000,64'b1100110000000000000000000000000000000000000000000000000000000000,64'b1110111000000000000000000000000000000000000000000000000000000000,64'b0111011000000000000000000000000000000000000000000000000000000100,64'b1111101100000000000000000000000000000000000000000000000000000000,64'b1111101110000000000000000000001000000000000000000000000000000000,64'b0100111111000000000000000000011110000000000000100000000000000000,64'b0011001111000000000000000000001010000000000000100000000000000000,64'b0000001101100000000000000000000111000000000000000000000000000000,64'b0000000100000000000000000001110000000000000001000000000000000000,64'b0000000000000000000000000000110000000100000001100000000000000000,64'b0000000000000000000000000000110111000010000111100000000000000000,64'b0000000000000000000000000000111101111110000000111000000000000000,64'b0000000000000000000000000011111100000111100000010000000000000000,64'b0000000000000000000000000011011100000001100000100000000000000000,64'b0000000000000000000000000001101110000000110000000000000000000000,64'b0000000000000000000000000000010001100000011111100000000000000000,64'b0000000000000000000000000000011001000000011110111000010000000000,64'b0000000000000000000001000000100000000000000111000110000000000000,64'b0000000000000000000011000000000000000000011011111111111000000000,64'b0000000000000000000001101110001111000000011000111111110000000000,64'b0000000000000000000000011000110011110000001001111001111100000000,64'b0000000000000000000011110110001000110000000001111111101100000000,64'b0000000000000000000001100000000110111001100001010000101000000000,64'b0000000000000000000000100110000111110000100000011101110000000000,64'b0000000000000000000000000010000111110001100011111111111100000000,64'b0000000000000000000000011010000011010000011110101000011111110000,64'b0000000000000000000000001110000011010110111100000001111111101000,64'b0000000000000000000000010110000101100110110000000001010011101000,64'b0000000000000000000000001100000000110010011000000001101101000000,64'b0000000000000000000000000000000000010010001000000011111111110000,64'b0000000000000000000000000000000000011000010000000010111110100000,64'b0000000000000000000000000000000000001100011010000010110000000000,64'b0000000000000000000000000000000000001100001110000010100000000000,64'b0000000000000000000000000000000000000010000110000010110000000000,64'b0000000000000000000000000000000000000011000110000100100000000000,64'b0000000000000000000000000000000000000011000010000100100000000000,64'b0000000000000000000000000000000000000001100011100101010000000000,64'b0000000000000000000000000000000000000001100010000110010000000000,64'b0000000000000000000000000000000000000000110001000100010000000000,64'b0000000000000000000000000000000000000000011101000100100000000000,64'b0000000000000000000000000000000000000000001100010101000000000000,64'b0000000000000000000000000000000000000000000100111011000000000000,64'b0000000000000000000000000000000000000000000100010100010000000000,64'b0000000000000000000000000000000000000000000110011011010000000000,64'b0000000000000000000000000000000000000000000110010111000000000000,64'b0000000000000000000000000000000000000000000110010111000000000000,64'b0000000000000000000000000000000000000000000110111010000000000000,64'b0000000000000000000000000000000000000000010111111010000000000000,64'b0000000000000000000000000000000000000000000011110110000000000000,64'b0000000000000000000000000000000000000000100000000110000000000000,64'b0000000000000000000000000000000000000000000011000010000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000100011100000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000010000000000000000000000000,64'b0000000000000000000000000000000000000010000000000000000000000000,64'b0000000000000000000000000000000000000010000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000100000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[93] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000111110000000000000,64'b0000000000000000000000000000000000000000011111111111000000000000,64'b0000000000000000000000000000000000000000000000000000010000000000,64'b0000000000000000000000000000000000000000011100000000010000000000,64'b0000000000000000000000000000000000000000000000000000011000000000,64'b0000000000000000000000000000000000000000000000000000001110000000,64'b0000000000000000000000000000000000000000001000000000000011100000,64'b0000000000000000000000000000000000000000000000000000000000110000,64'b0000000000000000000000000000000000000000000000000000000000001100,64'b0000000000000000000000000000000001111000000000000000000000000000,64'b0000000000000000000000000000001100000000000000000000000000000000,64'b0000000000000000000000000000000111111111000000000000000001000000,64'b0000000000000000000000000001111111111111110000000000000001100000,64'b0000000000000000000000000000111110000000000000000000000001100000,64'b0000000000000000000000000000000000000000000000000000000001100000,64'b0000000000000000000000110000000000000000000000000000000001101100,64'b0000000000000000000000111000000000000000000000001000000001110110,64'b0000000000000000000000100000000000000000000100000000000001100100,64'b0000000000000000000000000000000000000000000110000000000001100000,64'b0000000000000011000000000000000000000000000100000000000001100000,64'b0000000000000000000000000000000000000000000000000000000001110000,64'b1111111111111110000000000000000000000000000000000000000000100000,64'b0000000000000000000000000000000000000000000000000000000000100000,64'b1100000000000000000000000000000000000000000000000000000001100000,64'b0000000000000000000000000000000000000000000000000000000001100000,64'b0000000000000000001000000000000000000000000000000000000001000000,64'b1111111111111111000000000000000000000000000000000000000001000000,64'b1111111111111111111100000000111111000000000000000000000000000001,64'b0000000000000000000000000000001000000000000000000000000001110000,64'b0000000000000000000000000000111111000000000000000000010000111110,64'b0000000000000000000000000000000000000000111000000000000000000000,64'b0000000000000000000000000011111111111111111110000000000000000000,64'b0000000000000000000000000000011110000000000000000000000000000000,64'b0000010000000111111111000000000000000000000000000011111000000001,64'b1100111111100000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000010,64'b0000000000000000000000000000000000000000000000000111000001110001,64'b0000000000000000000000000000000000000000000000000000111111111000,64'b0000000000000000000000000000000000000000000000000000000000000111,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000111,64'b0000000000000000000000000000000000000000000000000000000000000011,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000011,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[94] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000010000000000000000000,64'b0000000000000000000000000000000000000000000001100000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b1000000000000000000000000000000000000000000000000000000000000000,64'b1111100000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111110000000000000000000000000000000000000000000000000000000000,64'b1111111000000000000000000000000000000000000000000000000000000000,64'b1000011100000000000000000000000000000000000000000000000000000000,64'b1000011100000000000000000000000000000000000000000000000000000000,64'b1010111100000000000000000000111110000000000000000000000000000000,64'b1100111111000000000000000000111100000000000000000000000000000000,64'b0010001111100000000000000001100100000000100000000000000000000000,64'b0011011111111000000000000011100111110001110000000000000000000000,64'b0011101101111100000000111110011111111110000000000000000000000000,64'b0000111111011100000010000011111111111101100000000000000000000000,64'b0001111111110000000000011111111100011111100000000000000000000000,64'b0000111111111000000100111110000000001000000001000000000000000000,64'b0000011111110000000001111000000000000000000000000000000000000000,64'b0000000000000000000111100000000000000000000000000000000000000000,64'b0000000000000000001111000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000001111100000000000000000,64'b0000000000000000100000000000000000000000001111100000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000001111000000000000000000,64'b0000000000000000000000000000000000000000111100000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000100000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000001100000000000000000000000000000000000000000,64'b0000000000000000000000100000000000000000000000000000000000000000,64'b0000000000000000000000011000000000000000000000000000000000000000,64'b0000000000000000000000111110000000000000000000000000000000000000,64'b0000000000000000000001111110000000000000000000000000000000000000,64'b0000000000000001111111111100001000000000000000000000000000000000,64'b0000000000000000000001111100001110000000000000000000000000000000,64'b0000000000000000000111111100000000000000000000000000000000000000,64'b0000000000000000000111110000000000000000000000000000000000000000,64'b0000000000000000011000000000000000000000000000000000000000000000,64'b0000000000000000111100000000000000000000000000000000000000000000,64'b0000000000000000011100000000000000000000000000000000000000000000,64'b0000000000000000110011000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000001000000000001110000000000000000000000000000000,64'b0000000000000000000000000000000111000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000001000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[95] = {64'b0000000000000000000000000000000000000000000001110010000110001000,64'b0000000000000000000000000000000000000000000000111100000110001111,64'b0000000000000000000000000000000000000000000000011111111110111001,64'b0000000000000000000000000000000000000000000000000011111110000000,64'b0000000000000000000000000000000000000000000000000000011110011000,64'b0000000000000000000000000000000000000000000000000000001111000011,64'b0000000000000000000000000000000000000000000000000000000011100001,64'b0000000000000000000000000000000000000000000000000000000000011000,64'b0000000000000000000000000000000000000000000000000000000000011000,64'b0000000000000000000000000000000000010000000000000000000000000111,64'b0000000000000000000000000000001111111111110000000000000000000000,64'b0000000000000000000000000000111111111111110000000000000000000000,64'b0000000000000000000000000000111110011111110000000000000000000000,64'b0000000000000000000000000000011111100111100000000000000000000000,64'b0011000000000000000000000000001111101100000000000000000000000000,64'b0000000000000000000000000111110011001110000000000000000000000000,64'b0000000000000000000000111111111110111110000000000000000000000000,64'b0000000000000000000001111100011111111110000000000000000000000000,64'b0000000000000000000001110100101111110000000000000000000000000000,64'b0000000000000000000111100000011101111100000000000000000000000000,64'b0000000000000000000111000000000000011100000000000000000000000000,64'b0000000000000000000110000000000000011100000000000000000000000000,64'b0000000000000000000110000000000000011110000000000000000000001111,64'b0000000000000000000110000000000001101111110000000000000000011111,64'b0000000000000000000111000000000111111111000000000000000000111111,64'b0000000000000000000111100000000001111111000000000000000000111111,64'b0000000000000000000111000000000111011110000110000000000001111001,64'b0000000000000000000111001111100000011000000100000000000000010011,64'b0000000000000000000111110001000010001100000110000000011111111111,64'b0000000000000000000111000000000000001100000110000001111111111001,64'b0000000000000000000111000000000100001100000110000011111111000000,64'b0000000000000000000011100100000101001100000110000011111111000000,64'b0000000000000000000011110110000100000111111100000011110000000000,64'b0000000000000000000001111011000011000101111110000011110000000111,64'b0000000000000000000000111101001111111111111100000000111110000000,64'b0000000000000000000000111000001010001111111110000111111110000000,64'b0000000000000000000000111000011001111111111000001111111110000000,64'b0000000000000000000000111111100010111100000000111111100000000000,64'b0000000000000000000000111000000000011100000001111011000000000000,64'b0000000000000000000000110000000010111000000001111000000000000000,64'b0000000000000000000001110001000100111000000001100100110000000000,64'b0000000000000000000001110001100111111000000001100101000000101111,64'b0000000000000000000001110001000111111000000011100001011111111110,64'b0000000000000000000001110000000011100000000010111111111111111111,64'b0000000000000000000001110000000011100000000001111111111100000001,64'b0000000000000000000001110000001011100000000000000011111110000000,64'b0000000000000000000001110000001111100000000000000000000110000000,64'b0000000000000000000001110000001111000000000000000000000100000000,64'b0000000000000000000001110100000011000000000000000000000000000000,64'b0000000000000000000001110101000011100000000000000000000000000111,64'b0000000000000000000001110100000111000000000000000000001100011100,64'b0000000000000000000011110101111111111100000000000000000110111111,64'b0000000000000000000001101111111111111100000000000000000111001111,64'b0000000000000000000000111111111110111100000000000000000011000111,64'b0000000000000000000000111111001111111111111110000000000011100100,64'b0000000000000000000000000010011111111001110000000000000011100001,64'b0000000000000000000000000011111111111111111100000000000011110010,64'b0000000000000000000000000000000000000000000000000000000001110000,64'b0000000000000000000000000000000000000000000000000000000001111110,64'b0000000000000000000000000000000000000000000000000000000001111010,64'b0000000000000000000000000000000000000000000000000000000000111110,64'b0000000000000000000000000000000000000000000000000000000000111111,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000101111111110000000000000000000000000000000000000000011111111};
assign input_o[96] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000010000100000000000000000000000000,64'b0000000000000000000000000000000010000100000000000000000000000000,64'b0000000000000000000000000000010010001100000000000000000000000000,64'b1111000001110000000000000000010010001100000000000000000000000000,64'b1000000001111000000000000000010010011100000000000000000000000000,64'b0000000000001000000000000000010110011100100000000000000000000000,64'b0000000000000000000000000000010010011100100000000000000000000000,64'b0000000000000000000000000000000010000110010000000000000000000000,64'b0000000111111111000000000000000010000100000000000000000000000000,64'b0000011111111111000000000000000010000100000000000000000000000000,64'b0000000111110000000000000000000010000100000000000000000000000000,64'b0000000000001111000000000000000010000100000000000000000000000000,64'b0000111111111111100000000000000010000100000000000000000000000000,64'b0000000000000000000111000000000010000100000000000000000000000000,64'b0000000000000000000011111000000010000000000000000000000000000000,64'b0000000000000000000000111000000000000000000000000000000000000000,64'b0000000000000000000000000000001100000000000000000000000000000000,64'b1111100000000000000000000000011111000000000000000000000000000000,64'b0000000000000000000000000000000000000000100000000000000000000000,64'b0000000000000000000000000000100000000011111000000000000000000000,64'b0000000000000000000000000011110000000000100000000000000000000000,64'b0000000000000000000000000011110000000000000000000000000000000000,64'b0000000000011111000000000001110000011000000000000000000000000000,64'b0000000000000000000000000001110000010000000000000000000000000000,64'b0000000000000000000000001001110000000000000000000000000000000000,64'b0000000000000000000000001110001111010000000000000000000000000110,64'b0000000000000000000000000110001000010000000000000000000000000000,64'b0000000000000000000000000111111000010000000000000000011111110000,64'b0000000000000000000000000111000001000000000000000000111111111110,64'b0000000000000000000000000111001001000000000000000011000000000000,64'b0000000000000000000000000111001111100000000000000011000011111111,64'b0000000000000000000000000111011100000000000000000000111111111111,64'b0000000000000000000000000111101000000000000011100000011111111000,64'b0000000000000000000000000011101000000000000000000000000000000000,64'b0000000000000000000000000011101000000000000000000000000000000011,64'b0000000000000000000000000001101000000000000000000000000000011111,64'b0000000000000000000000000011111100000011111100000000000000010000,64'b0000000000000000000111111111101110000000000000000000000000011111,64'b0000000000000000000100111101101110000000000000000000000000000000,64'b0000111111111000000110110001101110000000000000000000000000000000,64'b0000111111110000000111111001111100000000000000000000000000000000,64'b0000000000000000000000011101111001000000000000000000000000000000,64'b0000000000000000011000000000111000000000000000000000000000000000,64'b0000000000000000000000000000111100000000000000000000000000000000,64'b0000000000000000000000000000001111000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000001111111,64'b0000000000000000000000000000000000000000000000000000000000000001,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000111100000001100000000000,64'b0000000000000000000000100000000000000000000111100111111111111110,64'b0000011100111111111110000000000000000000000001111111000000000011,64'b0000000000000111100001111000000000000000000000111111111100000000,64'b0000000000000000000001000000000001000000000000001111111111000000,64'b0000000000000000000000000000111111111000000000000001101111110000,64'b0000000000000000000000000000011111111111000000000000000011111000,64'b0000000000000000000000000111110000000111000000000000000000000000,64'b0000000000000000000000000011111111110001111100000000000000000000,64'b0000000000000000000000000000011111111111000000000000000000000000,64'b1000000000000000000000000000000000111111111000000000000000000000,64'b0000000000000000000000000000000000000001100000000000000000000000};
assign input_o[97] = {64'b1110000000000000000000000000000000000000000000000000001100000000,64'b1110000000000000000000000000000000000000000000000000000100000000,64'b1110000111000000000000000000000000000000000000000000000000000000,64'b1110000010000000000000000000000000000000000000000000000000000000,64'b1110011100000000000000000000000000000000000000000000000100000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000111110,64'b1110000000000000000000000000000010000000000000000000000000001111,64'b1110000000000000000000000000000000000000000000000000000000000011,64'b1110000000000000000000000000000000000000000000000000000000000100,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1111000110000000000000000000000000000000000000000000000000000000,64'b1110000110000000000000000000000000000000011100000000000000000000,64'b1110000000000000000000000000000000000000000100000000000000000000,64'b1111000000000000000000000000000000000000000011000000000000000000,64'b1111000000000000000000000000000000000000000011111110000000000000,64'b1111000000000000000000000000000000000000000000000010011000000000,64'b1111000000000000011000000000000000000000000000000000111110000000,64'b1111000000000001111100000000000000000000000000011000011111110000,64'b1111000000000000001101000000000000000000000000000000000000011000,64'b1111000000000000001100000000000000000000000000000000000000001111,64'b1111000000000000001100000000000000000000000000000000001000000011,64'b1111000000000000000000000000000000000000000001100010000000000000,64'b1111000000000000000000111000000000000000000000111100000000000000,64'b1111000000000000000000111111111111110000001100110000000000000000,64'b1111000000000000000001000001110001111000001010001100000000000000,64'b1111000000000000000000000000000000000000000000100000000000000000,64'b1111000000000000000000000000000000000000000000100000000000000000,64'b1111000000000000000000000000000000000000010001000000000000000000,64'b1111000000000000000000000000000000000111110000000000000000000000,64'b1111000000000000000000000000000000000000010000000000000000000000,64'b1111000000000000000000000000000000000000000000100010000000000000,64'b1111000000000000000000000000000000000000001111011110000000000000,64'b1111000000000000000000000000000011111000000111111111000000000000,64'b1111000000000000000000000000000000000000000101111111000000000000,64'b1111000000000000000000000000100000111111000011100011000000000000,64'b1111000000000000000000000000100000011000000001110011000000000000,64'b1111000000011000000000000000000000111111100011110110000000000000,64'b1111001111111100000000000000000001111111100001111100000000000000,64'b1111111111111110001110110000111111111110000001001110000000000000,64'b1111000000000011111111000001110111111100000000000000000000000000,64'b1110000000000000000000000000010111111110000000000000000000000000,64'b1110000000000000000000010001101011111110010000000000000000000000,64'b1110000000000000000000111100000001101000000000000000000000000000,64'b0111111000000000000000111110111110101000000000000000000000000000,64'b1111100000000000011110001111111011111100000000000010000000000000,64'b1110000000000000000000000111111111111111111100000000000000000000,64'b1110000000000000000000000000011111111111111100000000000000000000,64'b1110000000000000000000000000000011111111110100000000000000001111,64'b1110000000000000000000000000000000001111111000000000000000000000,64'b1110000000000000000000000000000000000001111100000000000000000000,64'b1110000000000000000000000000000000000000000011100000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000,64'b1110000000000000000000000000000000000000000000000000000000000000};
assign input_o[98] = {64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000010000000000000000000000000000000000000000000000,64'b0000000000000000010000000000000000000000000000000000000000000000,64'b0000000000000000010011000000000000000000000000000000000000000000,64'b0000000000000000111111111111000100000000000000000000000000000000,64'b0000000000000000110011110000000000000000000000000000000000000000,64'b0000000000000000011111111110000000000000000000000000000000000000,64'b0000000000000000001111111110000000000000000000000000000000000000,64'b0000000000000000000000011100000000000000000000000000000000000000,64'b0000000000000000000000000111100000010111111000000000000000000000,64'b0000000000000000000000000011100000010011111000000000000000000000,64'b0000000000000000000000000111110111111101111000000000000000000000,64'b0000000000000000000000000110111101111111101110000000000000000000,64'b0000000000000000000000000011111111111111101111100000000000000000,64'b0000000000000000000000001111101111001111110001111100000000000000,64'b0000000000000000000000010000000011001000111111111110000000000000,64'b0000000000000000000000001100000011000000001111111110000000000000,64'b0000000000000000000000000110000001100111000111111110000000000000,64'b0000000000000000000000000010000001101111000011111110000000000000,64'b0000000000000000111100001010000001111111100001111011100000000000,64'b0000000000000010100110000011000000011101111000000001110000000000,64'b0000000000000110001011100011000000001111111000000011000000000000,64'b0000000000000011111101111111000000001110101000000000000000000000,64'b0000000000000001111111111100000000001111101000000000000000000000,64'b0000000000000000000111111100000000000001101000000000000000000000,64'b0000000000000000000001111000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000111100000000000000000000000,64'b0000000000000000000000000000000000000001110000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000010000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000010000000000000000000000000,64'b0000000000000000000000000000000000001000000000000000000000000000,64'b0000000000000000000000000000000000001000000000000000000000000000,64'b0000000000000000000000000000000000000111110000000000000000000000,64'b0000000000000000000000000001111000000000110000000000000000000000,64'b0000000000000000000000000000110000000110000000000000000000000000,64'b0000000000000000000000000000110000000000000000000000000000000000,64'b0000000000000000000000000000100000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000001100000000000000000000000000,64'b0000000000000000000000000000000000111000000000000000000000000000,64'b0000000000000000000000000000000001111000000000000000000000000000,64'b0000000000000000000000000000000000111000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000,64'b0000000000000000000000000000000000000000000000000000000000000000};
assign input_o[99] = {64'b0000000000000000000000000000000000000011110000000010000000100000,64'b0000000000000000000000000000000000000011111100000010000001111000,64'b0000000000000000000000000000000000000001111100000000000000101000,64'b0000000000000000000000000000000000000000110111000000000100011000,64'b0000000000000000000000000000000000000000110011000000010100001110,64'b0000000000000000000000000000000000000000110011000000010111100000,64'b0000000000000000000000000000000000000000011010100000000111110000,64'b0000000000000000000000000000000000000000011000111100000110100000,64'b0000000000000000000000000000000000000000110000111110000011000000,64'b0000000000000000000000000000000000000011110000000111000010000000,64'b0000000000000000000000000000000000000011100000001111100010000000,64'b0000000000000000000000000000000000000111111110000001100100000000,64'b0000000000000000000000000000000000000111000000000011101000000000,64'b0000000000000000000000000000000000000111000000000011011111110000,64'b0000000000000000000000000000000000000111000000000010111111000000,64'b0000000000000000000000000000000000000111000000000001110000000000,64'b0000000000000000000000000000000000001110000000000000100000000000,64'b0000000000000000000000000000000000001110000000000000000000000000,64'b0000000000000000000000000000000000001011000000000000000000000000,64'b0000000000000000000000000000000000001011000000001000000000000000,64'b0000000000000000000000000000000000001011010000111110000000000000,64'b0000000000000000000000000000000000001011010001111111100000000000,64'b0000000000000000000000000000000000001101100001110111000000000000,64'b0000000000000000000000000000000000000101100001101111100000000000,64'b0000000000000000000000000000000000000111100011101111111100000000,64'b0000000000000000000000000000000000000111011010011001111100000000,64'b0000000000000000000000000000000000001111100000011111101100000000,64'b0000000000000000000000000000000000011111000000111010110100000000,64'b0000000000000000000000000000000000011111000000000000111100000000,64'b0000000000000000000000000000000001111111110000000011000100000000,64'b0000000000000000000000000000000111001000000000001001100100000000,64'b0000000000000000000000000011111100011000000000000000111100000000,64'b0000000000000000000000000111111111110000000000000000011100000000,64'b0000000000000000000000001100000111100000000000000000000000000000,64'b0000000000000000000000011100000000000000000000000000000000000000,64'b0000000000000000000000110000011000000000000000000000000000000000,64'b0000000000000000001010100000110000000000000000000000000000000011,64'b0000000000000000011110100000000000000000000000000000000000000111,64'b0000000000000000111100001100000000000000000000000000001111111110,64'b0000000000000011100110001000000000000000000000000000001111111110,64'b0000000000000011001000100000000000000000000000000000001111000000,64'b0000000000000000011000000000000000000000000000000000001100000000,64'b0000000000000000000000000000000000000000000000100100011000000000,64'b1111111111111111111111111111111111111111111111111111111000000000,64'b1111111111111111111111111111111110011111111111111110011000000000,64'b1111111111111111111111111111111111111111111111101111011000000000,64'b1111111111111011111101101111111101111111111111111101110000000000,64'b1111111111111111111111111111111111111111111110111111110000000000,64'b1111111111111011111111111110111111111111011011111111100000000000,64'b1111111111111111111111111111111111111111111111111111100000000000,64'b1111111111111111111111111111111111111111111111111111100000000000,64'b1111111111111111111111111111111111111111111111111111000000001000,64'b0011000001111111011000011111000000010111111111100110000000000000,64'b0000011111100010000111100000000000001111111111001100000000000110,64'b1100011111101111000000000010000000111100101111011000000000000001,64'b0000001111001101100000000001000101110000011111010000000000000011,64'b0000000000001100001000000100000001010000010010100000000000000000,64'b0000000000001100000001111110000011000000000011100000000000000000,64'b0000000000001101000011111100000011000000001111100000000000000000,64'b0000000000110111000111101100010110000000001101100000000000000000,64'b0000000000000011000110001100011110000000000111100000000000000000,64'b0000000000001010001100001100001110000000000011000000000000000000,64'b0000000000001010001100001100101110000000000000000000000000000000,64'b0000000000001010001100001001001110000000000000000000000000000000};
endmodule
