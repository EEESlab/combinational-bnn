/* Module: data
 * Author: Manuele Rusci - manuele.rusci@unibo.it
 * Description: BNN net32 model stimulus.
 */


module data
(
	output logic [99:0][31:0][31:0] input_o
);
assign input_o[0] = {32'b00000000000000000000000000000000,32'b00000000000000000111011100000000,32'b00000000000000000101000000000000,32'b00000000000000000100111000000000,32'b00000000000000000011001100000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000111110001000000000,32'b00000000000011111111111100000000,32'b00000000000110111111101000000000,32'b00000000110001111011100000000000,32'b00000000110001101111000000000000,32'b00000000000000000110000000000000,32'b00000000000000000000110000000000,32'b00000000000000001010100000000000,32'b00000000000000000110100000000000,32'b00000000000000000010100010000000,32'b00000000000000000000100000000000,32'b00000000000000000111100001100110,32'b00000000000000001111111000000000,32'b00000000000000000110111000100100,32'b00000110000000000101110001000000,32'b00000111000000001011101111111100,32'b00000000001111111110010101111111,32'b00000000111111111111011111010110,32'b10000000000000001010100111111111,32'b00000000000000011111111110011110,32'b00000000000000011111100111111110,32'b00000000000000111001111110110110,32'b00001111111110001111011001111111,32'b00000111111111111000000111111111};
assign input_o[1] = {32'b00000000000000000000000000000000,32'b00000000000000000000111111000001,32'b00000000000000000000110111000111,32'b00000000000000000000110111000011,32'b00000000000000000000011110110011,32'b00000000000000000000001110011110,32'b00000000000000000000000000100001,32'b00000011000000000000000000000001,32'b00000011111001000000001100011111,32'b00000000000000000000000001111111,32'b11111110001111000001111111100000,32'b00000000011000011111110000000000,32'b00000000011000111111110000000000,32'b00001000111111101111110000000000,32'b00001011111000111011110000000000,32'b11111001111000111011110000000000,32'b11001001110000111011110000000000,32'b11101000110000011011000000000000,32'b11101111000000011111000000000000,32'b10011110100000011111000000000000,32'b00101000000000111110000000000000,32'b10111000000000111110000000000001,32'b00000000000000111100000000000111,32'b10000011000000101000000000011111,32'b00000000000001000000000011111011,32'b00000000000000000000001111011100,32'b00000000000000011001111111111000,32'b00000000000000000111101110000000,32'b00000000000000111100000000000000,32'b00000000000111100010000000000000,32'b00000000011110111000000000000000,32'b00000011110111000000000000000000};
assign input_o[2] = {32'b01110000000000000000000000000000,32'b01110000000000000000000000000000,32'b00100000000000000000000000000000,32'b00010000000000000000000000011111,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b10000000000000000000000000000000,32'b00000000000000010000000000000000,32'b11000000000111110000000000000000,32'b11100000000111111000000010000000,32'b11100000000111001110111111111000,32'b10000000000001101111011011110011,32'b00000000000001110111001100111000,32'b00000000000000110110000000000000,32'b11011100000000110111000000111111,32'b01111100000000011111000111111111,32'b11111100000000001000011111110011,32'b11110000001100011111111011000110,32'b01100000011111111100001111000000,32'b11000111111110011111100000000000,32'b00001111100111000001000000000000,32'b00001111110000000000000000000000,32'b10111110000000000000000000000000,32'b11100110000000000000000000000000,32'b11101110000000000000000000000000,32'b11011100000000000000000000000000};
assign input_o[3] = {32'b00000000000000000000000000001100,32'b00000000000000000000011111111011,32'b00000000000000000000000011111111,32'b00000000000000000000000000000000,32'b00100000000000000000000000111111,32'b11000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00011000000000000000000000000000,32'b00001110000000000000000000000000,32'b00000001100111111110010000000000,32'b00111111000011100000000000000100,32'b00000000000000001110000000000000,32'b00011111100000010000000000000000,32'b00000000000000001101000000000000,32'b00000000000001110110000000000000,32'b00000000000000001011000000000000,32'b00000000000000000010000000000000,32'b00000000000001111110011110000000,32'b00000000000011111100000000000000,32'b00000000000011111110000000000000,32'b00000111000011111111000000000000,32'b00000011111111111111100000000000,32'b00000000000111111111100000000000,32'b00000111001111001111100000000000,32'b00000000111111000011100000000000,32'b00000000011111001111100000000000,32'b00000000011011000000111100000000,32'b00000000000000110000001111000000,32'b10000000000000111111111110000000,32'b11000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[4] = {32'b00000000010000000000000000000000,32'b00000000001100000010000000000000,32'b00000000000000000000000000000000,32'b00000000000000101100001110000000,32'b00000000000000111001000100000000,32'b00000000111111100000001010000000,32'b00000000111111110000010000000000,32'b00000000010011100000000001000000,32'b00000000001111111111111101011000,32'b00000000000000000011111100010000,32'b00000000000000000000111110000000,32'b00000000001110000001000000001000,32'b00000000111100000011110000000100,32'b00000001011100000011100000000000,32'b00000111110100000010100000000000,32'b00000111100000000001100000000000,32'b10000111000000001110010000000000,32'b11111111011111111110000000000000,32'b11111111111111111110000000001111,32'b00000000010001111110000000000000,32'b00000000011011110110000000000000,32'b00000000011011111110000000000000,32'b00000000011011110010000000000111,32'b00000000001011111110000000011111,32'b00000000001011011110000000011111,32'b00000000001101111111000000111000,32'b00000000000111011110000000011110,32'b00000000000110001010000000001110,32'b00000000000011111000000000111111,32'b00000000000001100000000000010101,32'b00000000000000000000000000110100,32'b00000000000000000000000000111100};
assign input_o[5] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000011100000000000000000,32'b00000000000111110000000000000000,32'b00000000000001000000000000000000,32'b00000000000011111100000000000000,32'b00000000001110111100000000000000,32'b00000000000111011100000000000000,32'b00000000111111011110000000000000,32'b00000011101100010111100000000000,32'b00000110001100101111100000000000,32'b00000110001111111111010000000000,32'b00001100000101111111101100000000,32'b00001100100010111110011100000000,32'b00001110000010011100000011000000,32'b00001110011101100000010001100000,32'b00000110011100100000000001110000,32'b00001111001100010000000001110000,32'b00000111000000000000000001100000,32'b00000010011000111000001011100000,32'b00000010011001110000001111000000,32'b00000011110101111000001100000000,32'b00000001111001111000001100000000,32'b00000000011111111000011000000000,32'b00000000000000011000011000000000,32'b00000000000000001110110000000000,32'b00000000000000000100110000000000,32'b00000000000000001110110000000000,32'b00000000000000001100110000000000};
assign input_o[6] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000110000000000,32'b00000000000000000001100000000000,32'b00000000000000111101110000000000,32'b00000000000001111111111110000000,32'b00000000000011111111111111000000,32'b00000000000011111111111111000000,32'b00000000001111111001101111000000,32'b00000000001110111001100111000000,32'b00000000011111110011101111000000,32'b00000000011110110111111110000000,32'b00000000010110111101101110000000,32'b00000000001110011111111000000000,32'b00000000001100001111111000000000,32'b00000000001001010011110000000000,32'b00000000001101100111110000000000,32'b00000000011111100110000000000000,32'b00000000011111111110000000000000,32'b00000000011111111100000000000000,32'b00000000011111111000000000000000,32'b00000000110111111000000000000000,32'b00000001111110110000000000000000,32'b00000000111101100000000000000000,32'b00000000000001000000000000000000,32'b00000000000011000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[7] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000001000000000000000000000000,32'b00000001000000000000000000000000,32'b00000000001110000000000000000000,32'b00000000000000100000000000000000,32'b00000000011111110000000000000000,32'b00000010110011110000000000000000,32'b00000000101111000000000000000000,32'b00000000010011111000000000000000,32'b00000000011111111000000000000000,32'b00000000011111111000000000000000,32'b00000000000111111000000000000000,32'b00000000000011110000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00010000000000000000000000000000,32'b00010000000000000000000000000000,32'b00010000000000000000000000000000,32'b00001000000000000000000000000000,32'b00001000000000000000000000000000,32'b00001001000000000000000000000000,32'b00000001000000000000000000000000,32'b00000101000000000000000000000000};
assign input_o[8] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000001101100000111100,32'b00000000000000011100100000111000,32'b00000000000000001100100000111000,32'b00000000000000001000100000000000,32'b00000000000000001000000011111000,32'b00000000000000000000001111011011,32'b00000000000000000000110101110011,32'b00000000000000000011110001100001,32'b00000000000001111111100100011011,32'b00000000000001111111111000000000,32'b00000000000011111111100110000000,32'b00000000000011111111000000001000,32'b00000000000011101100000000011000,32'b00000000000111111100000000100110,32'b00000000000101010100000001001111,32'b00000000000101010000000000011111,32'b00000000000000000000000000111111,32'b00000000000000001000000001111111,32'b00000000000000000000000011111111,32'b00000000000000000000000001111011,32'b00000000000000000000000001111110,32'b00000000000000000000000011111110,32'b00000000000000000000000011111111,32'b00000000000000000000001111111010};
assign input_o[9] = {32'b00000110000000000000011000000000,32'b00000110000000000011111000000000,32'b10000111000000001111111000000000,32'b11111111000000000011111111100000,32'b11111111000000000001110111111000,32'b11111101000000000000000111101000,32'b00100101100000000000000000000100,32'b00001111111110010000000000000011,32'b00000111001111100000000000000000,32'b00000111110100010100000000000000,32'b00000001111111110100011111000000,32'b00000001101111111111111111000000,32'b00000000001111110000011111000000,32'b00000000000110000001010000000000,32'b00000000000110001100111111100000,32'b00000000000111111111111011100000,32'b00000000000110011111011110110000,32'b00000000000110110110110111100000,32'b00000000000011000000111000001001,32'b00000000000001111000001111001000,32'b00000000000001101000011010000011,32'b00000000000011111111111110000000,32'b00000000000011111000011111000000,32'b00000000000001101000011000000000,32'b00000000000011111111111001111000,32'b00000000000000111111101111111000,32'b00000000000001111111000000111100,32'b00000000000000000000000000011100,32'b00000000000000000000000000000000,32'b00000000000000000000000000011110,32'b00000000000000000000000000000111,32'b00000000000000000000000000010000};
assign input_o[10] = {32'b01100000000000000000000110100100,32'b00100000000000000000000110100100,32'b00000000000000000000000001111111,32'b00100000000000000000000001111100,32'b00100000000000000000000000001110,32'b00100000000111100000000000000111,32'b00000000000111110000000000000110,32'b00000000000111110000000000000011,32'b01000000000011001000000000000111,32'b00000000111111111111000000000011,32'b00000001111001111111100000000100,32'b01000001100000000101100000000000,32'b01000001101000000011100000011100,32'b01000001111100000111110000011100,32'b01000001111100001111110000010100,32'b00000000111100001111110000011111,32'b10000000101100001010110000001111,32'b10000000100100000010111000000110,32'b10000000011110111110101100000110,32'b00000000000111111111111010000011,32'b00000000000110111010011000000011,32'b00000000000111101011010000000000,32'b00000000000010101110000000000000,32'b00000000000010101110000000000000,32'b00000000000001100110000000000000,32'b00000000000001110011000000000000,32'b00000000000000101011000000000001,32'b00000000000000000111000000000000,32'b00000000000000000110000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[11] = {32'b00000000000000000000000000011010,32'b00000000000000000000000000011101,32'b00000000000000000000000000001110,32'b00000000000000000000000111101001,32'b00000000000000000000000101100011,32'b00000000000000000000000011001100,32'b00000000000000000000000000000000,32'b00000000000000000000011000000000,32'b00000000000000000000000000000000,32'b00000000000110000000000000000000,32'b00000000000000000001000000000000,32'b11111000000000011111000000000011,32'b10001111110000001101000000000000,32'b00011000001000111001000000000000,32'b00000000010101111111111111000000,32'b00000000001001100001110000111111,32'b00000000000101000000110100011000,32'b00000000110011000000110011111111,32'b00000000010111000000011110000011,32'b00000000010011110011110000000000,32'b00000000000000111011000000000000,32'b00000000000001111111101001000111,32'b00000000001001111110000011111111,32'b00000000001000011111111111111111,32'b00000000000010111110000000000001,32'b11000000000000100100000001110000,32'b01110000000000011100000000000000,32'b11001110000000000000000000000000,32'b00000111100000000000000000000000,32'b00001100110000000000000000000000,32'b00000011101111000000000000000000,32'b00000000111011110000000000000000};
assign input_o[12] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000001010000000000000000000,32'b00000000111111111110000000000000,32'b00000001111111111110000000000000,32'b00000000001000000111000000000000,32'b00011000000000000000100000000000,32'b00011000000001000000000000000000,32'b11100000000000000000000000000000,32'b10111111100000000000000000000000,32'b00000000111000000101100000000000,32'b00000000001000000000111000000000,32'b00001110000100000000110110000000,32'b00100000000000000000001111010001,32'b00000000000111010000000000000000,32'b00000000000001110000011111000000,32'b01110000000000000000000101100000,32'b11110011111100000000000000000000,32'b00000001110111110000000000000000,32'b00000000000111000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[13] = {32'b00000000000000000000000000000000,32'b00000000000000000011100000000000,32'b00000000000000000000100000000000,32'b00000000000000000001000000000000,32'b00000000000000000001110000000000,32'b00000000000000000001110000000000,32'b00000000111111000001111000000000,32'b00000000011101111111011000000000,32'b00000000011111111000111000000000,32'b00000000001100001111100000000000,32'b00000000001000000001000000000000,32'b00000000000000000001000000000000,32'b00000000001000000000110000000000,32'b00000000000101110000010000000000,32'b00000000000011000000000000000000,32'b00000000000000000000110110000000,32'b00000000000000100001111001110000,32'b00000000000001101111111100111100,32'b00000000000000111111111100000100,32'b00000000000001110111111100111100,32'b00000000000001110011111110111000,32'b00000000000000111111111111000000,32'b01100000000000111110111110000000,32'b01111111100000101110111110000000,32'b11111111110000100100011110000000,32'b01111000111111111100010110000000,32'b00111000111100011110011110000000,32'b00011111111001111111111000000000,32'b00111110101000000100000000000001,32'b11111101111110000000000000001111,32'b11110111101010000000000000011101,32'b11111111111011000001010011100110};
assign input_o[14] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000011100000000,32'b00000000001111100000001000000000,32'b00000000111011110000000100000000,32'b00000000101010100000000100000000,32'b00000000011001100010001100000000,32'b00000001111000111111000100000000,32'b00000111110011110000100000000000,32'b00000110111111110111100000000000,32'b00000110100000000001100000000000,32'b10000111111100000001100000000000,32'b00000101101000010001100000000000,32'b00001100011100011000110000000110,32'b11110111100000111000011000000100,32'b00000011111110000000011000000000,32'b00000001111110001110011000000000,32'b00000000000111001111001100000000,32'b00000000000011001101101100000010,32'b00000000000001100110111100000010,32'b00000000000000100110111100000000,32'b00000000000000110111110110000000,32'b00000000000000011011011110000000,32'b00000000000000011011011110000000,32'b00000000000000011111001111000000,32'b00000000000000001111001010000000,32'b00000000000000000111000110000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[15] = {32'b00000000000000000000000000000000,32'b00000011111000000000000000000000,32'b01000000000000000000000000111111,32'b11011000011111110000000000000001,32'b11100000000000000000000000000000,32'b11000000000000000000000000000001,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000010000000000000000000,32'b10000000001010000000000000000000,32'b10000000001000000001000000000000,32'b00000000000000000001000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00011111101000000000000000000000,32'b00000011100000000000000000000000,32'b01111000011000000000000000000000,32'b00111111001000000000000000000000,32'b10000001111000000000000000000000,32'b11111110001110000000000000000000,32'b00000001111111111100000000000000,32'b00000000000001011100000000010000,32'b00000000000000011100000000010000,32'b00000000000000001100000000000000,32'b00000000000000001000000000000100,32'b00000000000000000000000000000010,32'b00000000000000000000000000000001,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[16] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000001111001111111111000,32'b00000000000011111011111101111100,32'b00000000000111111011000000000000,32'b10000000000000000001111000000000,32'b10000011111000000001001100011000,32'b10111011110000000000001011000110,32'b00001110100000000001100001111111,32'b00000111110000000000000001111111,32'b00000111011100000000000111000001,32'b00000110010000000000001111000000,32'b00000111000100000000001110000010,32'b00000011000100000000000011111110,32'b11010011000010110000000011110000,32'b11100011000001100111100000001100,32'b01100010000000010000000111111101,32'b00000001110000001100000000000000,32'b00000000000000001100000000000011,32'b00000000000000000110000000000000,32'b00000000000000000001000000000000,32'b00000000000000000001000000000000,32'b00000000000000000001001100000000,32'b00000000000000000001001100000000,32'b00000000000000000001101100000000,32'b00000000000000000000111100000000,32'b00000000000000000000011000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[17] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000001111100000000000000000,32'b00000000011101111000000000000000,32'b00000000001111111000000000000000,32'b00000000000111111000000000000000,32'b00000000000011111011000000000000,32'b00000000001110001110100000000000,32'b00000001001111111111100000000000,32'b10011110011111111111100000000000,32'b10011011111110001111100000000000,32'b10000000111000000000011100000000,32'b00000000011110000000001011000000,32'b00000000001100000000000001100000,32'b00000000011100000000000011011111,32'b00000000011011000000000001111111,32'b00000011111111001010000000111111,32'b11110111111111101111111110111111,32'b11110011111000111100111110011100,32'b11110000101111111101111111110100,32'b00000000101111001110101110010001,32'b00000000011111111110100111111011,32'b00000000111111110000100001110111,32'b00011111011100000000000011111110,32'b11110111100000000000011111111000,32'b11111000000000000001111111110000,32'b10000000000000000000011110000000,32'b00000000000000000000010000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[18] = {32'b10000000000010000000000100100000,32'b10000000000000100000000011011000,32'b10000000000000111100110001100000,32'b10000000000000011110111100100000,32'b10000000000000000011110111111000,32'b10000001111111000111101001101000,32'b11110001111101100111101000111100,32'b11101111100000010111100000111100,32'b10001101110000011111100000111100,32'b10000111100000001111000000011000,32'b10000010000000000111100000000000,32'b10000010000000000100010000000000,32'b10000110000000000100000000000010,32'b10001110000000000101110000001001,32'b10001110000000000111000000001000,32'b10001010000000000011000000000000,32'b11101010000000000011000000111100,32'b10001110000000000001101110000001,32'b10000110000000000000110000000000,32'b10000110000000000000011000110000,32'b10000110000000000000001110000000,32'b10000011100000000111111011100000,32'b10000001100000000111110000110000,32'b10000001111111110110111100110000,32'b10000001111111111011101111111000,32'b10000000111111111101100011110000,32'b10000000000100001101110000110000,32'b10000000000000000111010000000000,32'b10000000000000000011111100000000,32'b10000000000000000011001100000010,32'b10000000000000000001111000000000,32'b10000000000000000000110100000000};
assign input_o[19] = {32'b00000000110010100011000000000000,32'b00000000111001010011000000000000,32'b00000000011001111111000000000000,32'b00000000001111111111000000000000,32'b00000000000101111000000000000000,32'b00000000000110110000000000000000,32'b00001111100011010000000000000000,32'b00001101100000100000000000000000,32'b00000111101111100000000000000000,32'b00000111000100000000001010010000,32'b00000011100000000000000000000000,32'b00000000000011110000001111000000,32'b00000000000001101000000110110000,32'b00000000110000010100000001100000,32'b00000000010000001000000000000000,32'b00000001111000100000000000000000,32'b00000000110000001110000000000000,32'b10000000000100011111000000000000,32'b11100000000011111011000000000000,32'b00100000000011110000100000000000,32'b11100000000011100100110000000000,32'b10100000000001111000010000010100,32'b11100000000000011100011000000000,32'b11100000000000001001111100100000,32'b11100000000000000000000101011000,32'b10100000000000000000001011000110,32'b10100000000000000000001111000000,32'b01000000000000000000000111000000,32'b01000000000000000000000011000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000100000000000000010000};
assign input_o[20] = {32'b00000010000000000011010100111110,32'b00011010000000000001010100111111,32'b10001110100000001001110110111110,32'b00000000000000000001101100111100,32'b00000000000000000001101100111100,32'b00000000000000000001011100111100,32'b00000000000000100111111111111100,32'b00000000000010111111110111111011,32'b00000000001111110011110000111000,32'b10000000111110001111110000011100,32'b00000111110110010111101111101111,32'b01111111101111111110000011111110,32'b11111111011101111111111100000000,32'b10111011101111100101100000000000,32'b10101110111111110011000000000000,32'b01001100000110110011000000000000,32'b00011111110111110010000000000000,32'b00001001111111100011000000000000,32'b00001111011111100111000000000000,32'b00100000000110001111000000000000,32'b11110000001111111011000000000000,32'b00000000000111101110000000000000,32'b00000000000011111011000000000000,32'b00000000000001111011000000000000,32'b00000000000000100011000000000000,32'b00000000000000001011000000000000,32'b00000000000000000000000000000000,32'b00000000000000001110000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[21] = {32'b01100010110110000000000001100010,32'b11111111111011111111001110010010,32'b01111001001101111011111010010010,32'b11111110001111111111100111010010,32'b11110110000011110001100111101000,32'b00111111110011110000000000110000,32'b11111111000000100000000000000000,32'b11011110000000110000000011111100,32'b11110000000000000100000011111011,32'b01001000000000000100001011111111,32'b00000000000000011100000101111111,32'b10000000000000010100010010110111,32'b00000000000000010111111111110000,32'b00000000000000111111111111110000,32'b00000000000000111011111111010000,32'b00000000000001011111111110010010,32'b00000000000000111110111111000000,32'b00000000000000111110111111000000,32'b00000000000100111111011110000000,32'b00000000000001100111011000000000,32'b00000000000001001010011111110000,32'b00000000000000001010011011010000,32'b00000000000000000110000110110000,32'b00000000000000010110000111110000,32'b00000000000000010000000000000000,32'b00000000000000010000000000000000,32'b00000000000000010000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[22] = {32'b00000000000000000000000110000000,32'b00000110101111100011111110000000,32'b00000110111001111111111000000000,32'b00000100000011110000000000000000,32'b00000000000111000000000000000000,32'b00000000000000000000000000000000,32'b11111110000000000000000000000000,32'b11111000111110000001000000000000,32'b10000000100111100000000000000000,32'b00000000001011110110000000000000,32'b00000000001110111000000000000000,32'b00000000001000011000000000000000,32'b00000000001000001000000000000000,32'b00000000001000001000000000000000,32'b00000000001000000001000000000000,32'b00000000011100001000000000000000,32'b00000000010100001000000000000000,32'b00000000001110000000000000000000,32'b00000000011110001111100000000000,32'b00000000010111011111100000000000,32'b00000000001111111111100000000000,32'b00000000000000000111011000000001,32'b00000000000000010111101000001010,32'b00000000000000000010010111001000,32'b00000011110000000010010101000000,32'b00000000000000000001111100000000,32'b00101000000000000001101100000000,32'b00100000000000000010000000000000,32'b01000000000000000001100000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[23] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000110000000000000000,32'b00000000000111111000000000101000,32'b01111000000011111000000000000100,32'b11111000000000011110000000000000,32'b11000111011111001111000000000001,32'b10000011111111111111111000000000,32'b00000010110000000001111000000000,32'b00000000011000000001111100000000,32'b00000111111000000011101100000000,32'b00000011111000000001000100000000,32'b00000000001000000001100000000000,32'b00000000011000000001100000000000,32'b11111000011000000000110000000000,32'b00000000011000000000110000000000,32'b00101000011000000000110000000000,32'b00100000001001111000110000000000,32'b00000000001101101001110000000000,32'b00000000000110100001100000000000,32'b00000000000011010001100000000000,32'b00000000000001010001100000000000,32'b00000000000000110111100000000000,32'b01110000000000000111100000000000,32'b00000000000000000001100000000000,32'b00000000000000000000000000000000,32'b00000000000000000001000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[24] = {32'b00000000000000100000110000000010,32'b01000000111111000010100000011100,32'b00111111110111101111100000001101,32'b11111111111111111110000000011110,32'b10111111111000000000000000001111,32'b10011110000000000000000000000000,32'b11110000000000000000000000000011,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000001011111111000000,32'b00000000000000000011111111100001,32'b00000000000011000001111111000010,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000011100000000000000,32'b00000000000000100000000000000000,32'b00000000000000000100001111111111,32'b00000000000111100100000000000111,32'b00000000000011111100011111111111,32'b00000000001111111100000000000000,32'b00000000000001111101100000000011,32'b00000000000000111100000011111111,32'b00000000000000000000111111111111,32'b00000000000100011111111111111111,32'b00000000000111111111111111111111,32'b00000001111111111101111110000000,32'b01111111111111111100000000000000,32'b11110111111111110000000000000000};
assign input_o[25] = {32'b00000000000000000000000000000000,32'b00000000001000000000000000000000,32'b00000001011000000000000000000000,32'b00000011011000000000000000000000,32'b00000001111000000000000000000000,32'b00000001111000000000000000000000,32'b00000001111000000000000000000000,32'b00000000110000000000000000000000,32'b00000001111110000000000000000000,32'b00000001001000000000000000000000,32'b00000001001110111111111110000000,32'b00000000111110011111111110000000,32'b00000001111100001111111100000000,32'b01100001001100001000000000000000,32'b00000000000100011000000000000000,32'b00000000000110011011101000000000,32'b00000000000011111101111001111111,32'b11110000000100000111101000000000,32'b00000000000111110100011000000000,32'b00000000000111100100001000001001,32'b00000001110110000000100111111111,32'b00000000111101100001110111000000,32'b11111111111100000001011100000000,32'b11111111110010000010001110100000,32'b00000000000000011110001100000000,32'b00000000000000001110011110100000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000111,32'b00000000000000000000000011111100,32'b11000000000000000111111100011111};
assign input_o[26] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000001111100000000000000000000,32'b00000001111100000000000000000000,32'b00000001001100000000000011110000,32'b00000001001100000000000001111000,32'b00000001101100000000000000000000,32'b00000101000011000000000000000000,32'b11100011000011000000000000000000,32'b01100001000011000000000000000000,32'b00000001001011000000000000000000,32'b00000000111111100000000000000000,32'b00000000111011100000001011110011,32'b00000000011111100000001111111111,32'b00000000001111011101111100000000,32'b00000000001111101111100000000000,32'b01111111111111111111100000000000,32'b00111111000100100110111000000000,32'b11110000000111100011111000000000,32'b00000000000111100000111111000000,32'b00000000000011100000111110000000,32'b00000000000111110000000000000000,32'b00000000000010110000000000000000,32'b00000000000001011100000000000000,32'b00000000000000111110000000000000,32'b00000000000000010000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000011111};
assign input_o[27] = {32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10110011111110000000000000000000,32'b11110110000010000000000000000000,32'b11101100000001000000000000000000,32'b11110111000001000000000000000000,32'b11100101100000100000000000000000,32'b10011111001100100000000000000000,32'b10111101111000110000000000000000,32'b10010110100000011000000000000000,32'b10000110000000001100000000000000,32'b10110000000000000110000000000000,32'b10110100000000000011000000000000,32'b10011000000000000001100000000000,32'b10001110000000000000110000000000,32'b10000110101110100000010001000000,32'b10000011101001100000011111000000,32'b10000000111000111100111111100000,32'b11100000000000000100101111100000,32'b10110000000000000011100011110000,32'b11011000000000000111000010100000,32'b10001100000000000011000000000000,32'b10000100000000000001100000000000,32'b10000110000000000001000000000000,32'b10000010000000000000100000000000,32'b10000000000000000000000000000000,32'b10000100000000000000000000000000,32'b10000100000111000000000000000000};
assign input_o[28] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000111100000000000000000,32'b00000000001111110000000000000000,32'b00000000001111001100000000000000,32'b00000000001111110000000000000000,32'b00000000001111100000000000000000,32'b00000000000000000000000000000000,32'b00000000000001100000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000001000000000000000000,32'b00000000000000000000000000000000,32'b00000000000111100000000000000000,32'b00100111000100000000000000000000,32'b00111000000100101100000000000000,32'b11100000000100011110000000000000,32'b00000000000000001111110000000000,32'b00000000000001111111111000000000,32'b00000000000000001111111000000000,32'b00000000000000011111011000000000,32'b00000000000000111110011000000000,32'b00000000000000000100000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[29] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000111110000000000000000,32'b00000000011111111111000000000000,32'b00000111111111011011000000000000,32'b00000111111111111011110000000000,32'b00000101000011111010111000000000,32'b00000110000000111110011000000000,32'b00001101111001111111111000000000,32'b00001101111100010111110000000000,32'b00000111110110010011111000000000,32'b00000111111100000101111100000000,32'b00000010101100000011011000000000,32'b00000011110100000010000000000000,32'b00000011011000001001010000000000,32'b00000011001100000000110000000000,32'b00000011001100111000000000000000,32'b00000011000111110110000000000000,32'b00000011000111111111000000000000,32'b00000011000011111111000000000000,32'b00000011000000111111100000000000,32'b00000010000000001101110000000000,32'b00000011011111000000010000000000,32'b00000011111111101000001100000000,32'b00000001011011111100000110000000,32'b00000001111000001111100111100000,32'b00000000111000000011100001100000};
assign input_o[30] = {32'b10010000000000000000000000000000,32'b10110000000000000000000000000000,32'b01100000000000000000000000000000,32'b11000000000000000000000000000000,32'b11000000000000000000000000000000,32'b11000000000000000000000000000000,32'b00000000111011100000000000000000,32'b00000000111111110000000000000000,32'b00000000010011111000000000000000,32'b00000000011011011000000000000000,32'b00000001111111001000000000000000,32'b00000001100010001010000000000000,32'b00000001111010101101000000000000,32'b00000000111110000110000000000000,32'b00000000111110010101000000000000,32'b00000000011110001111100000000000,32'b00000000001111111111100000000000,32'b00000000000001111110000000000000,32'b00000000000011110110000000000000,32'b00000000000000111110000000000000,32'b00000000000001111010100000000000,32'b00000000000001111001010000000000,32'b00000000000001101001111000000000,32'b00000000000000110100111100000000,32'b00000000000000001100011110000000,32'b00000000000000000000001100000000,32'b00000000000000000000000110000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[31] = {32'b00000000000000000000000000000010,32'b00000000000000000000000000000010,32'b00000000000000000000000000000010,32'b00000000000000000000000000000010,32'b00000000000000000000000000000010,32'b00000000000000000000000000000010,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000010,32'b00000000000000000000000000000010,32'b00000000000000000000000000000010,32'b00000000000000000000000000000010,32'b00000000000000000000000000000000,32'b11100000000000110000000000000000,32'b00000000000000000000000000000000,32'b11110000000000111110000000000000,32'b00000100000000011110000000000000,32'b11111000000110111110000000000000,32'b11111111110011101110000000000000,32'b01111111011111111000000000000000,32'b11111111000000111000001000000000,32'b00011110011111100110001000111111,32'b11111111111111110110000010111111,32'b11111111111111100010001001111111,32'b11111111111111100010011000000000,32'b11111110111001001010010001111111,32'b11100111111001010010010000011010,32'b11111110011001010010010001100001,32'b11111111010001010110000011000000,32'b11111001010011000000000000101111,32'b00000001010000000000000000011111};
assign input_o[32] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000011110000000000000000,32'b00000000000011111100000000000000,32'b00000000000001110110011100000000,32'b00000000000010000011001000000000,32'b00000000000011111001100000000000,32'b00000000000001100001110000000000,32'b00000000000001111100111100010000,32'b00000000000001100000001111000000,32'b00000000000001111010111100011111,32'b01111110000001100101111000011101,32'b00111110000001111111100000000000,32'b00000000000001111111000000000000,32'b00000000000011111111100000000000,32'b00000000000010011111100000000000,32'b00000000000011111111100000000000,32'b00000000000001111101000000000000,32'b00000000000000111110100000000000,32'b00000000000000001100110000000000,32'b00000000000000001101110000000000,32'b00000000000000001011110000000000,32'b00000000000000001111100000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[33] = {32'b00000000000011000001000000000000,32'b11111111111111000000000111111111,32'b10000000000001111000001111101111,32'b11111111111111110000000000001111,32'b11111111111111111111111111111111,32'b00000000000000000111111111110001,32'b01100000001111111011111111110000,32'b00000000001111110000011111110000,32'b00100000000011111110011111110000,32'b00000000000011111110000000000000,32'b00000000000000110010000000000000,32'b00000000000111000110000000000000,32'b00000000100000011100000000000000,32'b00000000100000001101110000000000,32'b00000000000000000000000000000000,32'b00000000000000000000111000000000,32'b00000000000001000000000000000000,32'b00000000001111000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000001100000000000000,32'b00000000000000010100000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000011110000000000000,32'b00000000000000011101000000000000,32'b00000000000000000011000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[34] = {32'b11000000000000000010001011100010,32'b11111100110000100010101011010010,32'b00000100000000100011101001010000,32'b00000011010000000011101001010000,32'b01000111010000000011101001111001,32'b00000001010000000011000001111000,32'b00000001111000000001001101111001,32'b00000011111000000001001100011011,32'b00000001101000001111111100000010,32'b00011111111000001000101000000110,32'b00001001111100000011110111100000,32'b00000011111100000000001111100000,32'b01000111111100000000001111000000,32'b11001100110100000000001111000000,32'b00110011111110000000000111100000,32'b00000001111100100000001110111110,32'b00000011111101000101111111111111,32'b00011110001011111110111111111111,32'b01001011111111101110001111111000,32'b01111111111111111111000000000000,32'b00111111111111111111000000000000,32'b11111111000011101101100000000000,32'b00111111111110101111000000000000,32'b00111001111000100011111100000000,32'b11111111111111111111111000000001,32'b11111111100000000000000000001100,32'b11111100000000001111000000000000,32'b11000000000000000000001000000000,32'b00000000000000001111100000000000,32'b00000000000000110000000000000000,32'b00000000001000000000000000000000,32'b01111111000000000000000000000000};
assign input_o[35] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000011110000101,32'b00000000000000000000011111100111,32'b00000000011111010001111111101111,32'b00000001110011111001110001111111,32'b00000111111111010001111011110000,32'b00000001001111111111111011110000,32'b00001111111111110000111001110000,32'b11111111111011111110011100110000,32'b11100001110001110110011010110000,32'b00001111110001110000011111110000,32'b11111111010011110000000111110000,32'b00000100111010110000000111010000,32'b00000000011010001110000000001111,32'b00000000011110001000000000011111,32'b00000000000111111110010000001111,32'b00000000000000001111111000000000,32'b00000000000000000000010000000000,32'b10000000000000001111100000111100,32'b00000000000000000000010000111111,32'b00000000000000000110000000111111,32'b00000000000001111111111111111000,32'b00000000001100111111111111000000,32'b00000000000001110000000000000000};
assign input_o[36] = {32'b00000000000000000000000000111110,32'b00000000000000000000000000111110,32'b00000000000000000000000000111110,32'b00000000000000000000000000111110,32'b10000000000000000000000000111110,32'b11100000000000000000000000111110,32'b11111100000111110000000000111110,32'b11111100011111111000000000111110,32'b11110110011101101111000000111110,32'b00011110011111111111000000111110,32'b00011011011111111111100000111110,32'b00001111001111111111100000111110,32'b00000111100011111000110000111111,32'b00000111110011111110110000111110,32'b00000011110011111110111000111110,32'b10000011011001100000111000111111,32'b11001111111001100000111000111110,32'b11110110111100111000011000111110,32'b11100011101111111000111000111110,32'b10000001001111011001111000111110,32'b00000000111011111111111100111110,32'b00000000001111111111110000111110,32'b11111100000000101111100000111111,32'b11111111111111101111000000111111,32'b00001000000011101110000000111110,32'b11111111111111111110000000111111,32'b11111111111111110010000000111111,32'b00100000000011111000000000111110,32'b00000000000000111000000000111110,32'b00000000000000111000000000111110,32'b00000000000000111100000000111110,32'b00000000000000111100000000111110};
assign input_o[37] = {32'b00000000000000001100000000000000,32'b00000000000000000011111111111111,32'b00000000000000000000000111110011,32'b00000000000000000000000111111110,32'b00000000000000000000000111110011,32'b00000000000000000000000000001100,32'b00000000000000000000000000000011,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000011111100000000000,32'b00000000000001111110000000000000,32'b00000000000001111111100000000000,32'b00000000000011000000000000000000,32'b00000000000011000000000000000000,32'b00000000000111111100000000000000,32'b00001111111100111100000000000000,32'b01100000001111110000011101100000,32'b11000000001100011100000000000000,32'b11100000000111100000000000000000,32'b00000000000000000011110000000000,32'b11000000000000101000000000000000,32'b01110000000000000010000000000000,32'b00011100000000111000000000000000,32'b00000111001111111111111111111111,32'b00000111110000000000000000011111,32'b00000110111110000000000000000000,32'b00000011101111111111111111111111,32'b00000000011001111110000000000000,32'b00000000001100000000000000000000,32'b00000000000001110000000000000000};
assign input_o[38] = {32'b00000000000000000000011000000010,32'b00000000000000000000011111111110,32'b00000000000000000000011100001111,32'b00000000000000001110001110000010,32'b00000000000011111111111110000001,32'b00000000000010111010011011100011,32'b00000000011110110000001111101101,32'b10000000001101111001111101111111,32'b00000000001111111111111111110000,32'b00000000000001001000011110010000,32'b00000000000001000001111000000011,32'b00000000000010111111111111110111,32'b00000000000010010001010111101110,32'b00000000000000010100111100011111,32'b00000000000011001110001100000001,32'b00000000000001010000111100000011,32'b00000000000000011111111000000011,32'b00000000000000011101111110111000,32'b00000000001110111111100111101000,32'b00000000001001010011100111111000,32'b00000000000000111111100111111100,32'b00000000000000110110001111111100,32'b00000000000000110100111110011111,32'b00000000000000010011111111000100,32'b00000000000000001111111111111110,32'b00000000000000001110000011011111,32'b00000000000001110110111111111111,32'b00000000000001110011111111111100,32'b00000000000011110000000011111100,32'b00000000000011111111100000011100,32'b00000000000000000000000000001110,32'b00000000000000000000000000000111};
assign input_o[39] = {32'b11000000000000000000000000000000,32'b01111110000000111111100000000000,32'b10111111011111111111111111000000,32'b11111110111111111000011111000000,32'b00011111111111111111111111000000,32'b11110111001111011111111111000000,32'b11000111111111111111111111000000,32'b00001001111001111111111110000000,32'b00001111001011011000000000000000,32'b00001111000001111000000000000000,32'b00011111011111010000000000000000,32'b00011011111000000000000000000000,32'b00001111011010000111000000000000,32'b00000111011010000011100000000000,32'b00001111011010000001100000000000,32'b00111111110111000001110000000000,32'b00110001110000000001110000000000,32'b00111111111011100111110000000000,32'b00010001111111110110000000000000,32'b00011011000000110110000000000000,32'b00001111001111111110000000000000,32'b00000010111111110110000000000000,32'b00000000001111111100000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000110000000000000,32'b00000000000000000000000000000000,32'b00000011000000000000000000000000,32'b11110000011111111111111111100000,32'b00000000000111110111111000000000,32'b00000000000000111011011111100000,32'b00001110111111110010111111100000};
assign input_o[40] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000001100000000000000000000,32'b11001100010100000000000000000000,32'b11111101111111000000000000000000,32'b01111000011110000000000000000000,32'b01111110010011111110000000000000,32'b00000011100001001110000000000110,32'b11001110010001000111000000000100,32'b11111110011101101101100000000000,32'b01000001111111110001110000000000,32'b00011000000011000101110000000111,32'b00010110000000000000111000000000,32'b01110111000000000001111000000000,32'b11110011000000000001100000000000,32'b11101010100000000001100000000000,32'b11101111110000000001100000000000,32'b11011111111111110001110000000000,32'b11001100111101001101110000000000,32'b11111100000110010110110000000000,32'b11111111000011010110110000000000,32'b11111111110111110111111100000000,32'b00000000111011010111111111000000,32'b00000000000111111001111110000000,32'b00000000000010101100011111000000,32'b01000001000000110111010000000000,32'b00000000000000011101010000000000,32'b00000000000000001111000000000000,32'b00000000111100000000000000000000,32'b00000001000100000000100000000000,32'b00000010000000000000110000000000};
assign input_o[41] = {32'b00000000000000000000000000000000,32'b11100000000000000000000010000000,32'b11111000000000000110111111111000,32'b11100000000000000111001111111000,32'b11110000000000000110011111111000,32'b01010000000000000110001110000100,32'b11000000000000000010001111111110,32'b01001000000000000011110000011111,32'b11111000000000001111100001001111,32'b11111000000111111011100000000011,32'b10110000000111111110000000000000,32'b11110000110000000000000000011111,32'b11111000000001111111000000000111,32'b11111000000010000111100000000001,32'b11011001111111000001000000000011,32'b11011001101110011000000000000000,32'b01011011100010100000000000000000,32'b01011011100001100110000000000000,32'b00111000100001100110000000000000,32'b01110010000001111110000000000000,32'b11101111110001110110000000000000,32'b00110111110001101110000000000000,32'b00001111000000101110000000000000,32'b00001100000100111110000000000000,32'b00010110111100000000000000000000,32'b00000010100000000000000000000000,32'b00000111111000000000000000000000,32'b00000111110000000000000000000000,32'b00000000100000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[42] = {32'b00000000000000000000000000000000,32'b00000100011111110000011000000111,32'b00000100000000000000000001000000,32'b10000100000000000000000111011111,32'b00000011111111111110000000000000,32'b00000000000011100000000000000000,32'b10000001111111111100000000001111,32'b00000000000000000000000000000000,32'b00001000111101111100000000000111,32'b00001000011011111100000000000100,32'b01001100001011011111100111111111,32'b00111101101111011110101100000111,32'b00001101101100000010011111000000,32'b00101101101100000000000000000011,32'b00101101101010000000010000001111,32'b00101100101110000001010011000000,32'b10100100101000000000010111000000,32'b00000100100000000011011110000000,32'b00100100110000000000011111000000,32'b11000110011101110000000000000000,32'b10111001111111111111011000001000,32'b11111111011111100110000000111000,32'b00011111111001111110000000111000,32'b00001111101111111111111111010111,32'b00000001111111111101111111101001,32'b00000000001111111001001110111111,32'b00000000000000111001000000111010,32'b00000000000000101000001011101111,32'b00000000000000101000000111100111,32'b00000000000000111100000111111010,32'b00000000111111101100001111111110,32'b00000001000000011110001111101110};
assign input_o[43] = {32'b00000000000010000000000010000000,32'b00000000000000000000000010100000,32'b00000000000000000000000100000000,32'b00000000000000000000000100000000,32'b00000000000000000000000101000000,32'b00000000000000000000000100000000,32'b00000000000000000000000000000000,32'b00000000000000000000001100000000,32'b00000000000101000000000100000000,32'b00000000000000000000000100000000,32'b00000000001111100000000100000000,32'b00000000000101000000000000000000,32'b00000000000111000000000000000000,32'b00000000000001000000000000000000,32'b00000000000001000000000000000000,32'b00000000000011000010000000000000,32'b10000000000011111111110000000000,32'b11100000000011111011110000000000,32'b11100000000011110001110000000000,32'b01000000000011011100000101000000,32'b11000000000111111111110100000000,32'b01000000000011111111111110000000,32'b10000000000001111111110000000000,32'b00000000000001100110000000000000,32'b10000000000001110111000000000000,32'b00000000000000101100000000000000,32'b00000000000000111011100000000000,32'b00000000000000011000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[44] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000111111000000000000000,32'b10000000001111111111100000000000,32'b10000000001111111000100000000010,32'b10000000001110111111001100000000,32'b10000000001110011101010000000000,32'b01100000001111111110111111111111,32'b01111000000111111011000000000011,32'b11111111111111111111111111110000,32'b11110000000111111111110000000000,32'b11111100000111110111111110000000,32'b00000100000011110000110001000000,32'b00000100000011111100000001000000,32'b00000100000111111100000001000000,32'b00000100000011111100000000000000,32'b00000000000011110110000000000000,32'b00000000000011001110000000000000,32'b00000000000011000101111111100000,32'b11111110000001000111111111110000,32'b00000000000001000001111111110000,32'b00000000000000011110000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[45] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000001111,32'b00000000000000000000000000000000,32'b00000000000000000000111111111111,32'b00000000000000000001111111111111,32'b00000000000110000001111000000000,32'b00000000000000000011111000000010,32'b00000011000000000011110000000010,32'b00000111100000111110110000000010,32'b00000011000000111000100000000010,32'b11111100000000011000100000000110,32'b11000001100000011111000011000111,32'b01111100100000111111100010001110,32'b01110111100000111111100000001110,32'b00011100110000111001110000001110,32'b11111111111110111001110000001110,32'b11101111110001111011100000000000,32'b11101100111111111111100000000000,32'b11111110000011111111100000000000,32'b11111111010011111110000000000011,32'b11111100000111111000000000101111,32'b11011100000111111000000000111000,32'b11011100000110111000000000101000,32'b01011100001111101000000000010000,32'b11111100011111111000000000010000,32'b10011100001110000000000000000000,32'b00000000001100000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[46] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b11111101001000000101110000000000,32'b11111111111111111100000001100000,32'b11111111111111111111111111110000,32'b00000000000011101101111000000000,32'b00000000001111010001100000000000,32'b00100100011111111001100000000000,32'b00111110111010111100100000000000,32'b00000000110011111100010000000000,32'b00000000111101111111110000000000,32'b00000000111111101111110000000000,32'b00000000011111111111110000000000,32'b00000000000001100000000000000000,32'b00000000000000100011111000000000,32'b00000000000000111111110000000000,32'b00000000000000111111101000000000,32'b00000000000000101111111000000000,32'b00000000000001010111111000000000,32'b00000000000011011111111000000000,32'b00000000011110001110001000000000,32'b00000000000011000000000000000000,32'b00000000000111110000000000000000,32'b00000000000011000111111000000000,32'b00000000011111000000110000000000,32'b00000000001100000001110000000000,32'b00000000000000000000000000000000,32'b00000000000000000000011110000000};
assign input_o[47] = {32'b10000000000000000001000000001000,32'b11000000000000000000100000100100,32'b11000000000000000000111111110001,32'b11000000000000000000001111110001,32'b11000000000000000000000011100100,32'b11000000000000000000000001100111,32'b11011111000000000000000011110000,32'b10011100000000000000000000000001,32'b10111000111100000000000000000000,32'b11111110010110000000000000000000,32'b11111111000011000000000000000000,32'b11011101100001000000000000000000,32'b10000111110001100000000000000000,32'b10000101101100100000000000000000,32'b10110110111110110000000000000000,32'b10011001011111010000000000000000,32'b10110000100110110000000000000000,32'b11111011011011011111000000000000,32'b10001100001000111111010000000010,32'b10001100010000001111010000000000,32'b10000111111111111101111100000000,32'b10000111111111111001100000000000,32'b10000000001111111100110010000000,32'b10000000000000001111111100100000,32'b10000000000000000111101110100000,32'b10000000000000000011111111100000,32'b10000000000000000000111111000000,32'b10000000000000000000001100000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000000000000000000};
assign input_o[48] = {32'b00000010000000000000000000000000,32'b00000110000000000000010011111000,32'b00000000000001100000011111110011,32'b00000011100001100000010111000111,32'b00001000111110000111101100110111,32'b00000011110000001111111111111110,32'b00000000000000000111000111101110,32'b00000000000000011110000110100110,32'b00000011000011111110111111001110,32'b11101000111111101111111111111111,32'b11001101110111111100000011000010,32'b11011000111100000000000000000000,32'b11110011100000000000000000000000,32'b10110000000000000000000000000000,32'b00100000000000000000000000000000,32'b11111000000000000000000000000000,32'b00000000000000001100000000000011,32'b11000000000000010001100000000011,32'b11110000000000010010110000001111,32'b11110000000000000110010011111000,32'b11110000000010001111011110000111,32'b00100000001101101111110001111111,32'b00000000000010101101111111111011,32'b00000000000000011001110011111110,32'b00111111111111111111111111100000,32'b11111110001110001100010000000000,32'b10000011010011111011110000000000,32'b00000010010010011101111111000000,32'b00000000011010111100001110000010,32'b10000001010010011000001100001110,32'b00000010011111110010011100001000,32'b00000010001110110000000010000000};
assign input_o[49] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000001111111110000000000,32'b00000000000101111111110000000000,32'b00000000011111111111111100000000,32'b00000000010110000000001100000000,32'b00000011111100000000001100000000,32'b00000110111100000000000110000000,32'b00000110110110000000000100000000,32'b00001101111110000000011110000000,32'b00001101111110000000010110000000,32'b00111000001100000000010010000000,32'b00011000010100000000000010000000,32'b00110000011000000000010000000000,32'b00100111111001100001111100000000,32'b00011111111011100001110000000000,32'b00000111111110100011000000000000,32'b00000000111011100011100000000000,32'b00000000111111100110000000000000,32'b00000000101111000100000000000000,32'b00000000001101001100000000000000,32'b00000000000000101000000000000000,32'b00000000000000011000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[50] = {32'b00000000000000000000000000000000,32'b00000001000000001111111111111111,32'b00000101111111111101111111111111,32'b11000100001111111111111110000000,32'b11111111111100000000000000000000,32'b00000000111000000000000000000000,32'b00000001111100000000000000000000,32'b00000000111111100000000000000000,32'b00000000011110100000000000000000,32'b00000000000111110000000000000000,32'b00111000111001110000000000000000,32'b00111111001001010000000000000000,32'b11100000001000010000000000000000,32'b00000000001001111000011000010100,32'b00000000001011111000000000011111,32'b00000000001110111000001100101010,32'b00000000001101111000011111101110,32'b00000000001110101100001101001110,32'b00000000011111110110000000001100,32'b00000000011110011011000000001000,32'b00000000011110011101100000000000,32'b00000000010100000101111110000100,32'b00000000101111110111001110000000,32'b00011111111011000011011111110000,32'b11000000011000001100010111111111,32'b00000000001111001111111110000000,32'b00000000111111100000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[51] = {32'b11110000000000000000000000000000,32'b11110000000000000000000000000000,32'b11110000000000000000000000000000,32'b11110000000000000000000000000000,32'b11110000000000000001111000000001,32'b11110000000000011111111100000000,32'b11111110000000000111111111000011,32'b11111110000000000111111111111000,32'b11111100111111111101111111111000,32'b11111111111111111111000001111111,32'b11111111100011100000000000000111,32'b11110000000111000010000000000000,32'b11110000000000010000000000000000,32'b11110000000000000000000000000000,32'b11110000000000000000000000000000,32'b11110000000000000000000000000000,32'b11111111111111100000001100000000,32'b11111000000000000110001111000000,32'b11110001111111110001101111110000,32'b11101000011110001100111110000011,32'b11110000001110000100000000000011,32'b11110000000000000100000000000000,32'b11110000000001111100000000001000,32'b11110000000000000000000111111000,32'b11110000000000000000001110000000,32'b11110000000000000000111000000000,32'b11100000000000000011100000000000,32'b11110000000000001111000000000000,32'b11110010000000111101000000000000,32'b11110000000011110100000000000000,32'b11110000001110000000000000000000,32'b11110001111100000000000000000000};
assign input_o[52] = {32'b00100110000011010000000000000000,32'b00011111111101111111111000000000,32'b00000011100111000111111111100000,32'b00000000001111111110001111111111,32'b00000000000111001000111110111111,32'b00000000000011011111011111111101,32'b00000000111111111011111011110111,32'b00000111111111111111111000000111,32'b00000111111100011111111000000000,32'b00000011111111111111110000000000,32'b00000001111101111111110000000000,32'b00000000110000011111111010000000,32'b00000000011000111111111010000000,32'b00000000000001011111101101000000,32'b00000001111000111101000110100000,32'b00000000110110011111100011010011,32'b00000000011001110011110000101110,32'b00000000011010110011111000010111,32'b00000000001101111111011000001111,32'b00000000011111111111101110001110,32'b00000000010111101110111010001110,32'b00000000001011111101011111101110,32'b00000000000101001100001101111100,32'b10000000000000100001011111111100,32'b10000000000000000001111111111100,32'b01100000000000000001111111111000,32'b11001000000000000000111111111011,32'b00010010000000000000111111110001,32'b00000100011100000000010101110001,32'b00000000110001000000000011111000,32'b00000000000000011100000011111011,32'b00000000000000011000000011111010};
assign input_o[53] = {32'b11110000000000000000000000000000,32'b11111101000000000000000000000000,32'b11111110000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000001111110000000000,32'b00000000000000011100000010000111,32'b00000000000001111101111001101110,32'b00000000000011111110000000000001,32'b11110000001111111111111111111111,32'b11111111111111111111111111110010,32'b11000000001111111111000111000000,32'b11111111111111111111111110000000,32'b00000000001111111111000010000000,32'b11111111111011101111011110000000,32'b00000000100000111111000000000000,32'b00000011001111101000000010000000,32'b00000010000011011000000000000000,32'b00000000011111110000000000000000,32'b11111111111111110110000000000000,32'b00011111111111111110000000000000,32'b11111111111111100000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[54] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b11000000000000000000000000000000,32'b01000000000000000000000000000000,32'b10000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b01100000000000000000000000000000,32'b11100000000000000000000000000000,32'b11100000000000000000000000011111,32'b11100000000000000000000000011111,32'b11000000000010000001100011111111,32'b00000000000010101001111111100000,32'b00000001000001000001110000000000,32'b00000000000110001111110000000000,32'b00111111111110011111100000000000,32'b00011001111111110111100000000000,32'b11111111110101101111000000000000,32'b11011111111111011111000000000000,32'b00001111100011111111000000000000,32'b00001101100111111110000000000000,32'b00000101000111101111000000000000,32'b00001110000111111111000000000000,32'b00010010001111101111000000000000,32'b00001100000011011111000000000000,32'b00001110000011000111000000000000,32'b00000000000000011100000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000001111,32'b00000000000000000000000001111110,32'b00000000000000000000001111111111,32'b00000000000000000001111111111100};
assign input_o[55] = {32'b10101100000000000000000000000000,32'b11111100000000000000000000000000,32'b11111011100000000000000001000000,32'b11111000000000000000000001010000,32'b11111000000000001100000001010000,32'b11111000000000011100000001111000,32'b00111000011000011100000000111000,32'b00010100111100010111110000111000,32'b00000000111111001111110000000000,32'b00000000101111011111111100000000,32'b00000000000011111111011110000000,32'b00000000000001111110000100000000,32'b00000000000111110110001111010000,32'b00000000000100111111111100000000,32'b00000000000101111111101110100000,32'b00000000000101111011111111111111,32'b00000000000001001100111111110110,32'b11000000000000011000011010001111,32'b00000000000000001111110010000000,32'b00000000000011111111011011111110,32'b00000000000000001101011100110110,32'b00011111000000001111011111011100,32'b00001111111111100111101011010001,32'b00011111111111001010100110110110,32'b00000111110011111001100000001111,32'b00000011110001110011111000011111,32'b00000001111111110001101000000000,32'b00000000111110011110000000000000,32'b00011111111111111010000000000000,32'b00111111111000111110000000000000,32'b00111111011011111111000000000000,32'b01111010111111110111000000000011};
assign input_o[56] = {32'b00000000000000000000000000011100,32'b00000000000000000000000000000111,32'b00000000000000000000000000011101,32'b00000000000000000000001101111111,32'b00000000000000000000111110110001,32'b00000000000000000001111111110111,32'b00000000000000000011100011101111,32'b00000000000000000011000011111101,32'b00000000000000000011100111111100,32'b00000000000000000011101110001100,32'b00000000000000000011101100110110,32'b00000000000000001111111111111111,32'b00000000000000011011000001111111,32'b00000000000011110100100001110111,32'b00000000000110111111100000001111,32'b00000000001111111111000000000011,32'b00000000000111100000000000000011,32'b00000000001100000000000001110101,32'b00000111111110000000000001111000,32'b00011111111110000000000001111011,32'b00111111111110000000001011001111,32'b00101111001100000000000000011111,32'b00010000111000000000111001111111,32'b11111111111111111111001011111011,32'b11111111111111111101111111101111,32'b11111111111111111111111011011110,32'b11111111111111111111111111111100,32'b11111111111111111111111101111100,32'b00000011000001000001111000111101,32'b00000011000111000001111000001010,32'b00000010000011000000110100001010,32'b00000110001110000000010110011100};
assign input_o[57] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000011111000000,32'b01111111100000011111111111111111,32'b00000001111111110000001110011111,32'b00000011111100000000000000000001,32'b00000000110111111000000000000000,32'b00000000111011110000000000000000,32'b00001110000111100000000000000001,32'b00011000011110000000000000000011,32'b00000000010011111000000000000111,32'b00001000001011000000000011111110,32'b00000111001011000000000011110011,32'b00000000001101110000011111100001,32'b00000011100111000000111000000000,32'b00111111110011100111110000000000,32'b11111100111111010000111000000000,32'b10000011110011110011111100000000,32'b10000011010001110111111110000000,32'b11000001111000110111111110000001,32'b11000001101101111011011100000000,32'b11100000111010001101111110000000,32'b11100000011110000100011000000000,32'b11100000011110000011001110000000,32'b11110000001101111110101111000000,32'b11111000001111100011110110000000,32'b11111100000110110001111000000000,32'b01111100000011111000011110000000,32'b10111110000011111111100000000000,32'b11011010000001101110100000000000,32'b11101111000000111111100000000000};
assign input_o[58] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000011111100000000000000,32'b00000000000011111110000000000000,32'b11111100000001111110000000000000,32'b11111111100000111110000000000000,32'b01111001100000011100000000000000,32'b00000001100000000000000000000000,32'b00000011111100000000001100000000,32'b00000011111000000000110000000000,32'b00011110111000000000101000000000,32'b11111111111000000000101000000000,32'b00111001110000000000101100000111,32'b00000001010000000000011100011111,32'b00000001011000000001111100001111,32'b00000000101000000000111111110011,32'b00000011111000000000000111110000,32'b00000001111000000000000000010000,32'b00000001111000000000000001100000,32'b00000001011000000000000001100000,32'b00000011011000000000000000100000,32'b00000011110000000000000000000010,32'b00000011110000101000000000000000,32'b00000010100000000000000000000000,32'b00000110100000100000000000000000,32'b00000111100000000000000000000000,32'b00000111100000000000000000000000,32'b00001111000000000000000000000000};
assign input_o[59] = {32'b00000000000001000000000000000000,32'b00000100000001011100111111111000,32'b00000100000001001100111111111111,32'b00000100000001001111111110111111,32'b11111100000001001011111111111111,32'b00011100000000001111110000000000,32'b01111100100000001000000000000000,32'b11100000000000000000000000001111,32'b10001111100000001111111111111111,32'b00111111110000111111100011001000,32'b00000110000000000111100000000000,32'b00001110000000001111000000000000,32'b00000000000000000011000000000000,32'b00000000000001111111000000000000,32'b00000000000000111000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000010000000000000000,32'b00000000000000000000000000000001,32'b00000000000000000000000000000111,32'b00000000000000101000000011111110,32'b00000000011101111111111111100000,32'b11100001110001111111110000000000,32'b11111100011111110000000000000000,32'b11111111110000010000000000000000,32'b11111111100011111000000000000000,32'b10001000001111000000000000000000,32'b00000000000000110000000000000000,32'b00000000000000000011000000000000,32'b00000000000000000000001110000000};
assign input_o[60] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000010000,32'b00001101000000000000000000000000,32'b00000100000000000000000000000000,32'b00000100000000000000000000000000,32'b00000100000000000000000001100000,32'b00010101000000000000000000100000,32'b00000100000000000000000000000011,32'b00111100000011111111111111111100,32'b01101100000011110000111110000111,32'b11101011100001100110111010000000,32'b11011111100000101110000001111000,32'b01101111100000001110111111000000,32'b11100111110010001110100001000000,32'b01000110110000001110111000000000,32'b01100111100010001110100000000000,32'b11111111110011111110101001110000,32'b11100111100111011110011111110000,32'b11111111100001111110001100110000,32'b00011101100001101110001111110000,32'b11111111000001011110001111011000,32'b01110111000001110110001101011000,32'b11110101000000110110000100010000,32'b11100111000000010110000110010000,32'b00101100111000000100000000110000,32'b00001111000000000011111000100000,32'b11111111110000011110011000000000,32'b00000110000011110011111000000000,32'b00111000111101111110000000000000,32'b00011110011111100000000000000000,32'b11100111110000000000000000000000,32'b11111100000000000000000000000000};
assign input_o[61] = {32'b01101000000000000000000000000000,32'b01111000000000000000000000000000,32'b00111000000000000000000000000100,32'b11110110000011000000111000010100,32'b00000011110100011000010001101100,32'b01100101110101110000000010101100,32'b00000101110011011111100101110111,32'b00101100000000000000011101110000,32'b10111100001101111111110010000000,32'b00011111100011111111111111110001,32'b00000010011110111110111011111100,32'b00001111001111111111111101111100,32'b00000000111111101000011111111100,32'b00000000000010000011111011111000,32'b00000000000001101111011001111010,32'b00000000000000000000011111110111,32'b00000000000000111111111101101000,32'b11000000000001111111101111100000,32'b11000000010000111111101111101000,32'b10000000000001101111001111111101,32'b10100000000001111111001111111111,32'b00001000000001111011001111110000,32'b10111100000001000111000111101111,32'b11110111110000011110111111111110,32'b11011011110100001000001111111111,32'b11111101111010000011000011111111,32'b11000111111111111000010000000000,32'b00000000010111111110010000000000,32'b00000000001111111111100000000000,32'b00000000000011111111111100000000,32'b00000000000000000111011111000000,32'b00000000000000000111111111110000};
assign input_o[62] = {32'b00000000000000000000111010000000,32'b00000000000000111110011010000000,32'b00000000000000111110001110000000,32'b00000000000000111110000100000010,32'b00000000100000011110000010010000,32'b00000000100000011100000001111000,32'b00000000100000000000000000111111,32'b00000000000000010100000000111111,32'b00000001000001111100000000111111,32'b00000001000000111100000000000011,32'b00000001000011111111100000000011,32'b00000001000111101111110000001010,32'b00000000000110000010110001111000,32'b00000000001101000011111111111000,32'b00000000001101000011111110111000,32'b00000000001101001011111111111100,32'b00000000001111111011111111111000,32'b00000000001111110111111100011110,32'b00000000000111111011111000010100,32'b00000000000000111111100001111110,32'b00000000000000111011100001101110,32'b00000000000000111011100001111110,32'b00000000000000011001100000111110,32'b00000000100001100111100111101011,32'b00000000000000000111100000011100,32'b00000000000000001011111111111111,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[63] = {32'b00000000010000010000000000000000,32'b00000000000000010000000000000000,32'b00000000000000010000000000000111,32'b00000000000000010000000000010000,32'b00000000000000010000000000011111,32'b00000000000000010000000000111100,32'b00000000000000010000000000110000,32'b11100000000000010000000001110000,32'b11100001000000010000000011110011,32'b11100111101111010000000000110111,32'b11100111101011010000000000110110,32'b11100111101010011000000000110110,32'b11100010100000011000110000110111,32'b01100010100000001100000001111011,32'b11100010101000111100100001111111,32'b11100110000001111100110001111000,32'b11000001111011101100000001111011,32'b00000000000011111100111011111001,32'b01000110000001111110101001111011,32'b00011111111111111111111111111100,32'b11000111101111111000011101101111,32'b00011111111111111111000111111101,32'b00000000000000111000000111111111,32'b00000000000000000001000000000111,32'b00000000000000000000000000000000,32'b00000000000000001000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[64] = {32'b00000000000000000000000000000000,32'b01000111110000111111100000000111,32'b11100000110000000000100000000001,32'b00000000011000001111100000000001,32'b00000000010000000000000000000110,32'b00000000000111000000000000111111,32'b00000000111001111111100000001110,32'b00000000111111011111111000000011,32'b00000000000111111111100000001111,32'b11100001011111000011100000011111,32'b01111001110001111101000000010100,32'b01111000110011110110011111111110,32'b11111001000000000000000000001101,32'b10000111000000000000000000001101,32'b01111111100000000011000000001100,32'b11111111110111111110000000000100,32'b00000011111001111010000000000110,32'b01110011111101010010000000000011,32'b00000111011101010010000000000001,32'b00111111011101100010000000000000,32'b00101111111101100010000000000000,32'b11100111100001100110000000000000,32'b11101110000000100110000000000000,32'b11111110000000011111111111000000,32'b11111110000010001111111100000000,32'b10110100000001000011111111000000,32'b01110100111000100000000000000000,32'b00001011011101100000000000000000,32'b00001100111111100000000000000000,32'b11111111000000000000000000000000,32'b01111100100000000000000000000000,32'b11111111110000000000000000000000};
assign input_o[65] = {32'b00000000010111101101000101000000,32'b00000000001001101101111111111100,32'b00000000000001110101111111111001,32'b00000000100111111000000000011000,32'b00000000100000010000000001111111,32'b00000000100111111100000001111111,32'b00000001100111111000000001111011,32'b00000001000111111100000000000000,32'b00000001000011110000000000011100,32'b00000001000011111110000011111110,32'b00000000000001111110000011101100,32'b00000000000000000100000011111111,32'b00000000010111111111000001111000,32'b00000000010110000011000000111000,32'b00000000001100011001000001111000,32'b00000010100011111001110000111000,32'b00000000111110111101110000011000,32'b00000000111111101101110001100000,32'b00000000111110111101110000110000,32'b00000000011111110111100000000000,32'b00000000000001100000000000100000,32'b00000000100001100000000010000000,32'b00000000000001100000000011111110,32'b00000000000000100000000010111000,32'b00000000000000011111111111111110,32'b00000000000000000000000011111100,32'b00000000000000010110000001111111,32'b00000001000000000000000000000000,32'b00000001000000000000000000000000,32'b00000000000000000000000000000000,32'b00000010000000000000000000000000,32'b00000010000000000000000000000000};
assign input_o[66] = {32'b10000000010000000000100000000000,32'b10000000010000000000110000000000,32'b10000000011000000000011000000000,32'b10000000001101000000001110000000,32'b10000000000110000000000111100000,32'b10000000000011100000000001110000,32'b11000000000000111000000000011000,32'b11111000000000001111000000011100,32'b11011100000000000000100000000100,32'b11000110000000000000110000000111,32'b11000011100000000000001000000111,32'b11000001100000000000000111000010,32'b11000000100000000000000001110010,32'b11000001110000000000000000011011,32'b11000000110000000000000000001111,32'b11000000110000000000000000001111,32'b11000011100000000000000000001010,32'b11100001000000000000000000011010,32'b11011101111100100000000000000110,32'b11110111100111110000000000110011,32'b11011111100001111000000000000000,32'b11111111111100111111000100001100,32'b11111111111111011110111111000000,32'b11110011111111101111100000000000,32'b11000000000011111101110000000000,32'b11000000000000111111110110000000,32'b11000000000000001111101110000000,32'b11000000000000000011100110000000,32'b11000000000000000000000000000000,32'b11000000000000000000000000000000,32'b11000000000000000000000000000000,32'b11000000000000000000000000000000};
assign input_o[67] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000111110000000000000000000000,32'b00001000000000000000000000000000,32'b00011111110000000000000000000000,32'b00000000000000000000000000000000,32'b00001000000000000000000000000000,32'b00001000000000000000000000000000,32'b00000011110000000100000000000000,32'b00000000000000000100000000000011,32'b00000000000000111100000000000001,32'b00000000000000001100000000000001,32'b00000000000000000000000000000000,32'b00000000000000011100000000000000,32'b00000000000000000100000000000000,32'b00000000000000011111000000000000,32'b00000000000000001100000000000000,32'b00000000000000111100000000001111,32'b00000000000000000100000000011110,32'b00000000000000000100111110111111,32'b00000000000011111000111111111110,32'b00000000000011111111111111110000,32'b10000001111100111111000001111111,32'b11111111111000000000011111111100,32'b11111000000100111111111100000011,32'b00000111111100000000000000000000,32'b01111111111100000011100000000000,32'b11111000000000000000000000000000,32'b00000111100111000000000000111100};
assign input_o[68] = {32'b00010000000000000000000000001110,32'b01110000000000000000000001011111,32'b00000000000000000000000001011100,32'b00000000000000000000000001011100,32'b10100000000000000000110001011100,32'b10101000000000000000000000111100,32'b10101000000000000000000000111111,32'b00111000001110000011110000011111,32'b00111000001000000111111111101100,32'b00111100000100000111111110001111,32'b00110101001011110110011100111111,32'b00010101001101111011111111111111,32'b00011100000011100100011100011111,32'b00011110010000000001111111111100,32'b11011110000000011010111111100000,32'b11001100110011111100001000000000,32'b11000111111010111110000000000000,32'b01000001111001100000000000000000,32'b00000000000111011110000000000000,32'b11110011000010111110000000000000,32'b01010000111111011110000000000000,32'b01011111111111111110000000000000,32'b11110011111111100000000000000000,32'b11100000011111100000000000000000,32'b11111111100001100000000000000111,32'b11111111100111000010000000111111,32'b01111111111111100000000000110111,32'b00111111100000000000000001111111,32'b00000000000000000000000000001111,32'b00000000000000000000000010000000,32'b00000000000000001000000000000000,32'b00000000000001110000001110000000};
assign input_o[69] = {32'b00000011000000100111000000000000,32'b11111011011100101111111001100111,32'b10001011110011111110011001111000,32'b00111111111111111111011110000000,32'b11110001100111111101111000000000,32'b10011111111101110011100000000000,32'b00000010100101010000000000000000,32'b00000001101011110000000000000000,32'b11111111100100000000000001111111,32'b10001111111001110000000000000000,32'b10001111010000001110000000000000,32'b11100111110000010100000000000000,32'b11110000010000010000000000000000,32'b11000000000000010000000000000000,32'b11100000000000011110000000000000,32'b00000000100011111110000000000000,32'b00000000000111101110000110000000,32'b00000000001110001100000110000000,32'b00000000000011111100000000000000,32'b00000000000001111100000000000000,32'b00000000000111100000000000000000,32'b00000000000001111110000000100000,32'b00000000000000000000000000000000,32'b00000000000000100000000000100000,32'b00000000000000100000000000000000,32'b00000000000000011111000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[70] = {32'b00000000000000000000000000000000,32'b00000000000000000000011111111111,32'b00000000000000000000000000000000,32'b00000000000000000000000000000001,32'b00000000000000000000000000011100,32'b10000000000001111000000000000000,32'b11000000000001011000000000000000,32'b10000000000011111000000000000000,32'b10000000000011111000000000000000,32'b10000000011111100111100000000000,32'b00000000010000000111110000000000,32'b00000011110000000010111000000000,32'b11111001110000000000001100000000,32'b01101011111000000001111100000000,32'b01110100110000000001110000000000,32'b11010011100000000000110000000000,32'b11111111100000000000111100000000,32'b00011000011111000000110000000000,32'b00000000000100111000111000000000,32'b00000000010111111000110000000000,32'b00000000010010000000110000001111,32'b00000000011011000000110000111100,32'b00000000001111000000101111110000,32'b00000000000010000011111111111110,32'b00000000000110000010100001110000,32'b10000000000010000000111000000000,32'b10000000000111111110101000000000,32'b10111000000110011110111000000000,32'b11111011001100000011111000001011,32'b00001000001100011111110101111100,32'b00001100011011111111111111100000,32'b00000100000011111100111100000000};
assign input_o[71] = {32'b10000000000000000000000000000000,32'b10000100000000000000000000000000,32'b10000000000000000000000000000000,32'b10000000000000000100000000000000,32'b11000000000000000000000000000000,32'b10111110001100000000000000000000,32'b11111111000100100000000000000000,32'b10110010010010000100000000000000,32'b10110110100001100110000000000000,32'b10011110100000110000000000000000,32'b10001101100000011000000000000000,32'b10000000000000001000000000000000,32'b10011000110000000100000000000000,32'b10000000110000000110000000000000,32'b10000000010000000110000000000000,32'b10000000011000000011000000000000,32'b10000000001000000011110000000000,32'b10000000000000000000011000000000,32'b11100000000000000000011000000000,32'b10011000000001110000001000000000,32'b10000110000000011110000100010000,32'b11101110000000111011100000000000,32'b10000110000001100100111001000000,32'b10000011111101001110000111000000,32'b10000000001011000000000011100000,32'b10000000000111000000000111100000,32'b10000000001101101000000111100000,32'b10000000101111111000000011100000,32'b11110000111111111000000101110000,32'b11111111001100101000000000000000,32'b10111001101111010000000000000000,32'b11000111111111011100000000011100};
assign input_o[72] = {32'b00000000000000000000000000000000,32'b00000000000000000001100111111111,32'b00011111111000000000000000000000,32'b11111111000000111110010000000000,32'b00000000000011111100001000000000,32'b00000000000000000000000000000000,32'b01111000000000010000100000000000,32'b11111111100000000001111110000011,32'b11111111111111010011100000001110,32'b10000000000011110000010000000111,32'b11000000010001111110000000000000,32'b01111111100000100010000000000001,32'b00000000000011100011100000000000,32'b00000000000111100011000000000000,32'b00000000000101110001110000000000,32'b00000000000011110001110000100000,32'b00000000000010111111111111000011,32'b00000000000001111110111111111000,32'b00000000000111111111111111100111,32'b00000000000011111101000000001111,32'b00000000000001110101000001111000,32'b10000000000001110101000000000000,32'b00001111000000111111000000000000,32'b00100000000000111011100000000000,32'b10101111111000100101100000000000,32'b11100000000000001100011111100000,32'b00000111100000000000111111111111,32'b11000011111111111100001111000000,32'b10000000000000001111111111111111,32'b00000000000000000000000000000000,32'b11100000000000000011000000000000,32'b10100000000000000000000000000000};
assign input_o[73] = {32'b00000000001011000000000000000000,32'b11110000011111000111110000011110,32'b00111110000100011000000000000000,32'b11000000000000000001110000000000,32'b00000000011111000000000000000000,32'b00000000000011100000000000000000,32'b00000000000111001111110000000000,32'b11100000000011001011111000000000,32'b11100000100010110111011100000000,32'b10000000100010000000111000000000,32'b00000000100000000001111000000000,32'b11000000100000000000110000000000,32'b00000001100000000000110000000000,32'b00000001000000000000110000000000,32'b00000001000000000000110000000000,32'b01100001000100000000001100000000,32'b00011001001100000000000100000000,32'b01101001101000000000111100000000,32'b00000011001000000001110000000000,32'b11001011111110100000110000000000,32'b00110011111111110000010100000000,32'b00000000101111111100010100000000,32'b00000000011001011111111011000000,32'b00000001100000101101111000000000,32'b00000001110011111111111000000000,32'b00000001101111010111111000000000,32'b00000001011111110011100111111111,32'b00000001011101111111100000001100,32'b00110001000100111111111111111111,32'b00010011000111111111111111111111,32'b00001111111111111111101111111111,32'b00001100111111100000000000000000};
assign input_o[74] = {32'b00000000000000000000000001001110,32'b01000000000000000000000001011111,32'b00000000000000000000000001011100,32'b00000000000000000000000001011000,32'b00000000000000000001100001011100,32'b00100000000000000001110001011100,32'b00100000000000000000110001011111,32'b00101000000100100000000001001110,32'b00101000001001111100000000111111,32'b00111000001011111111101111111100,32'b00111100000001111111001000011111,32'b00010100001111111111111001111111,32'b00010100111111110011110111111111,32'b00011100011110000000111111111111,32'b00011100011110001111111111111100,32'b10011110001110111111110111100000,32'b10011100010111111111110000000000,32'b10001111101101111111110000000000,32'b10000000000111110010100000000000,32'b11000111111111111110100000000000,32'b10111111011011000011110000000000,32'b11110111111011010111110000000000,32'b11110111011111100101110000000000,32'b11111111111101111111110000000000,32'b11011111111111111000000000000000,32'b11010000000111110000000000000000,32'b11101111111111000000000000000000,32'b11111111111011000000000000111111,32'b11111111111111000000000000111111,32'b00111111111000000000000000011111,32'b00000000000001110000000000001111,32'b00000000000000000000000000000000};
assign input_o[75] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000001111100000000,32'b00000000000000000001111100000000,32'b00000000000000000000100110000000,32'b00000000000000000001110111000000,32'b00000000000000001111111011000000,32'b00000000000000011111011101011111,32'b00000000000000010111111111111110,32'b00000000000000010000111011111111,32'b00000000000000000001111111110101,32'b00000000000000000100111110000001,32'b00000000000000000000111000000000,32'b00000000000001111001111000000011,32'b00000000000001001111100000001111,32'b00000000000011101111110001111110,32'b00000000000111000001111011111100,32'b00000000001111100000111111100000,32'b00000000111110000010000000000000,32'b00000000001110010000010000000000,32'b00000000100110000000000000000000,32'b00000000100000000000000000000000,32'b00000000100000000000000000000000,32'b00000000000000000000000000000000,32'b00000001111000100000000000000000,32'b00000000000000011111000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[76] = {32'b00100000000000000000000100100000,32'b00101000000000000000000100100000,32'b00101000000000000000000001100000,32'b00101000000000000000000001100000,32'b00001000000000000000000001100000,32'b01100000000000000000000000100000,32'b01110011000000000000000001100000,32'b00010111000000000000100001100000,32'b11110011000001000000000000100000,32'b00110110000001001111000000100000,32'b11100010000001100111111111100000,32'b00000111110100110111110111100000,32'b11111111100000011011111000000000,32'b10010011110011110111111100100001,32'b00000001100111111111011100000100,32'b00001111110110000111111100001000,32'b00000000000000111011110000000000,32'b00000000000001111011110000000000,32'b00000000000001111011111111110111,32'b00000000000001111000111111111100,32'b00000000000001111101101000001111,32'b00000000000000101111111111110011,32'b00000000000000110000000000000001,32'b00000000000000011111111111110000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000011100000};
assign input_o[77] = {32'b11100000000111000000000000000000,32'b11100000000111000000000000000000,32'b11100000000111000000000000000000,32'b11110000000110000000000000000000,32'b01101000000011100111111111000000,32'b00111000000000000000000011111111,32'b11111100000010000001100000001100,32'b11111111110000100000000000000111,32'b11011111000011111001100000000100,32'b11001111111110000000000000000000,32'b11111111111111111111111100011000,32'b11101111000111111111111000011100,32'b11111000000001100000000000001000,32'b11100000011100110000000000000111,32'b11100000011111011100000000000100,32'b11100000011111001000000000000011,32'b11100000011111001000000000000000,32'b11110000000001001000000000000111,32'b11111111011000011110000000010000,32'b01111101111111111111111000111111,32'b11111111111110011111111111111111,32'b11111111101110111110111111111100,32'b11111111111100011001111100000001,32'b11111111001111111111111000000010,32'b01111110111111000000000000000001,32'b11100111111100100000000000000000,32'b11101111000000000111111100000000,32'b11100000000001111111111000000000,32'b11100000001111100011110000000000,32'b11100000001000001100000000000000,32'b11100000001110000000000000000000,32'b11100000000000000000000000000100};
assign input_o[78] = {32'b00000000000010000000001001001010,32'b00000000100010010100000011000111,32'b00000000000010010100000000000111,32'b11000000000010010000110010000111,32'b01000000000000001100110000000001,32'b01000000000000000111110000000000,32'b01000000000000000011010000001000,32'b01000000000000000001100000001000,32'b00000000000000000000110000000000,32'b10000000000000001100010000011000,32'b10000000000000111110000100000000,32'b10000000000000110111000110000000,32'b10100000000011100101000111111111,32'b00000000000011001111111111011110,32'b00000000000011011111101011000000,32'b00000000000011101111101111100100,32'b00000000000011110011000011100110,32'b00000000000001111111110011111111,32'b00000000000001110111100001111110,32'b00000000000000111111100000000010,32'b00000000000000111101000000000000,32'b00000000000000010011000001000000,32'b00000000000000010001000000000000,32'b00000000000000001111000000000000,32'b00000000000000000011000000011111,32'b10000000000000011100100000000000,32'b00000000000000000100000000011111,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[79] = {32'b00000001000000000000000000000000,32'b00000011000000000000000000000000,32'b11110001000000000000000000000000,32'b11100000000000000000000000000000,32'b00100001000000000000000000000000,32'b00100011110000000000000000000000,32'b11110001100000000000000000000100,32'b11111111100000010000011000010100,32'b01111111111110011100000000110110,32'b11001111000110011100011001010100,32'b10001001011110001111000001010110,32'b11111000110111111000001000110001,32'b01111000011111111000000100000100,32'b00000001101111111110000100000001,32'b00000011111111110110000010000010,32'b00000000101111111110000000000010,32'b00000000000111111010001010000010,32'b00000000111011111101001010000010,32'b00000000000101111100111001000010,32'b00000000000000111001101101100010,32'b00000000001111101111111100111010,32'b00000000000010100001100011001110,32'b00000000000000011111111111000010,32'b00000000000011101111111111110010,32'b00000000000001001111111111111001,32'b00000000000000010000001000000100,32'b00000000000000000000000000000000,32'b00010111000000000000000000000000,32'b00001111110000000000000000000000,32'b00000111011100000010000000000000,32'b00000001110111000000000000000000,32'b00000000011111110000000000000000};
assign input_o[80] = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000001110000000000,32'b00000000000000000000100000000000,32'b00000000000001100000111000000000,32'b00000000000011110000010000000000,32'b00011111110011111110011100110000,32'b00000000000001111111100010000001,32'b00111110000000011110000011111100,32'b00000000000000000000000000001111,32'b11100000000000000000000011111111,32'b00011111000000000000000011000000,32'b11110000000000000000111100000000,32'b00000000111101010111111100011110,32'b00000000011111111111001011111111,32'b00111111100111111111010000111111,32'b00000000000111111111000000011111,32'b11111111010000011111111111111111,32'b10111111110111111110001001100000,32'b11111111111111100100000001000000,32'b10000111111111100000000000000000,32'b01100000000001100000000000000001,32'b00000000000001000000111000000000,32'b00000000111111100001111000000111,32'b00000000000001100000011000000011,32'b00000000011000000000000000011111,32'b00000001110000000001001111111111,32'b00000000010111111111111111011111,32'b11111111110000001011111111111111,32'b11111010011111111111000000000000};
assign input_o[81] = {32'b00000000000000000000111010000010,32'b00000000000000000000110110011111,32'b00000000000000000000110001111111,32'b00000000000000000000111101000110,32'b00000000000000000000110101111110,32'b00000000000000000000110101000011,32'b00000000000000000001110101100010,32'b00000000000000000011000000100000,32'b00000000000000000011110000110000,32'b00000000000000000000110110110010,32'b00000000000000111100110111010001,32'b00000000000000111110100100110010,32'b00000000000000111110001011110010,32'b00000000000000110110011001110001,32'b00000000000000101110111010110000,32'b00000000000001101011111011111111,32'b00000000000001101011011111111111,32'b00000000000001101111111111111111,32'b00000000000001111111110111111111,32'b00000000000011011111000011111111,32'b00000000000011010011000000010011,32'b00000000000010111111000000000000,32'b00000000000000111111110000000000,32'b00000000000000001110111000000000,32'b00000000000000000111111000000000,32'b00000000000000000000010000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[82] = {32'b00000000000000000000000000000000,32'b00000001111000000000000001111111,32'b00000000001100000001110011111111,32'b01100000000000000000000011101111,32'b10000000000000000111000000000111,32'b10000000000000001010000000000000,32'b11111111001100111111000000000000,32'b10000000110001111110000000000000,32'b10101111100011111110000000000000,32'b11111111111111110110000000000000,32'b00000000011111011111010000000000,32'b00000000011111101111100000000000,32'b00000000111111100101000000011111,32'b00000000111011000111100000011111,32'b00000000111100000011000000000111,32'b00000010101110000011101111111111,32'b00000111001100001111110000001111,32'b10000111101110000111100000000000,32'b00000101111111111111100000000000,32'b00000001001111111100000000000000,32'b00000001111111011111000000011100,32'b00000001111111111000000111111000,32'b00000001111111110110000000011111,32'b00000000010111111100000000000000,32'b00000000000111100000000000000000,32'b00000000000011100000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[83] = {32'b00000000000000000000000000000000,32'b00000000000111100000000001111111,32'b00000000000000000000000011000000,32'b00000000000000000000011100000000,32'b11111000000000000000111100100111,32'b00000111000000000000011110100000,32'b00000000100000000000011110000000,32'b00000000000000000000000010000000,32'b11111111100000000000000100001111,32'b11111111100000000000000011111110,32'b11111111000000000000000001111000,32'b01111100000001111100000011111100,32'b11101010000001000000000001111000,32'b01101010000000011111000011111111,32'b01001010000000011010100101000000,32'b00001010000111100001100011000000,32'b11111110000111111100000000000011,32'b01100011001110111100000000000000,32'b11100010000011111100000000011110,32'b11101100000001001100000000000000,32'b11100100101000001000000000011111,32'b11100000001000000000000000010000,32'b00100000000000010000000000000000,32'b00011000000000000000000000111111,32'b00011000000000000000000000000000,32'b11001111000000000000000000000000,32'b11111100000000000000000000000000,32'b11111000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[84] = {32'b00010101001000000000000000000000,32'b11111111111111111110000011111111,32'b00010000000111111111011011110000,32'b11011111111111111110000001111110,32'b01111111111111111101111110000011,32'b11111111111111001011111111111111,32'b01100111111111111111000000000000,32'b01111111011110111111111111111111,32'b11111111111110011001111111011111,32'b11111110001110110000000000111111,32'b11111111111111111111011111100111,32'b11111111110110000010011111111100,32'b11111111101110011110000011111111,32'b00000000110111100010111111101000,32'b00000000001101111111111111111111,32'b00000110011001100010011111111101,32'b00000000000001100000000000111111,32'b00000110010000100000001111100111,32'b00000000110000100101101111110010,32'b00000000000000101101111001110111,32'b00000000000000100101111111111011,32'b00000000000000100100011111111011,32'b00000000000000000000000011111111,32'b11100000000000010000000000000001,32'b11100000000000000000011111000000,32'b01100000000000000011111111110000,32'b11111100000000000000000110000000,32'b11010011111111111111111110000000,32'b00001111111111111111011111100000,32'b11111111111111111111111111000110,32'b11111111000000000000001111111000,32'b11100000000000000000000000011111};
assign input_o[85] = {32'b00000000000000000000000000100000,32'b00000000111111110011111110011000,32'b00000000000000010000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000100000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000011111,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000001100000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00110000000000000000000000000000,32'b11110000000000001100000000000000,32'b00111110000000001100000000000000,32'b11111000000000010000000000000000,32'b00000000000000010000000000000000,32'b00000111100000000000111111111111,32'b00000011111000000011111111111111,32'b11111111110000000011111000000111,32'b11111001111000000000000000010000,32'b11111111111000000000000001100000,32'b11111111000000000000011100011111,32'b11000000000000000000000001111111,32'b00000000000000000000111111111100,32'b00000000110001111111111111001100,32'b00000000111111111110011111110000,32'b00111111111111111100100000000000};
assign input_o[86] = {32'b00000000000000000000110001100000,32'b00000000000000000000110001000000,32'b00001101110000000011100001000000,32'b11100001100110000000100010000000,32'b00000111111111110011100011000000,32'b00110111111111100011000010000000,32'b00000011100110000111000000000000,32'b00000011111101000010000100000000,32'b00000000110011111111000100000000,32'b00000001110001011111100000000000,32'b00000001100000110111100000000000,32'b00000011100000000011100000000000,32'b00000011000000000011000000000000,32'b00000001100000010011000000000000,32'b00000000110000000011000000000000,32'b00000111111111000001000000000000,32'b00000000100001000001100000000000,32'b00000100111111100000100000000000,32'b00000000110111000000110000000000,32'b00000000110000000001100000000000,32'b00000000111000111111100000000000,32'b00000000011111111101110000000000,32'b00000000110111000110111000000000,32'b00000000011001000001111000000000,32'b00000011111111001000110100000000,32'b00000111011101000000011010000000,32'b00000011000011101000000101110000,32'b00000000000011000000000011110000,32'b00001000001110100000000000000000,32'b00001110001000100000001111000000,32'b00001110010000000000001110000000,32'b00111001000001100000011010000000};
assign input_o[87] = {32'b11000000000000000000000000000000,32'b11000000000000000000000000000000,32'b11000000000000000000000000000000,32'b11000000000000000000000011100000,32'b11000000000000000000000100110000,32'b11000001100000000000000000000000,32'b11000111111000000000000000000000,32'b11000011111000000000000000001011,32'b11000011101111110000000000000111,32'b11000000101111111100000000000110,32'b11000001100000111110000000000111,32'b11000000100000001111000000111000,32'b11000001100000000011100110000000,32'b11000011110000100001100000001111,32'b11000001110000000011110000110000,32'b11000000111000000001101110000000,32'b11000000011111000000111000000000,32'b11000001011111000000111100000000,32'b11011111101111000011111110000000,32'b11000001111100110011011110000000,32'b11001110010100101111111110000000,32'b11110000000011110111111000000010,32'b11000000000000111111111100001110,32'b11000000000000011111111111000000,32'b11000000000000000111111111110001,32'b11000000000000000111111111000000,32'b11000000000001111001111111010000,32'b11000000001111000111111110100000,32'b11000000000000001000011110111000,32'b11111111000001110000000111111111,32'b11010000001110000000000000110110,32'b11000011111000000000000000011100};
assign input_o[88] = {32'b00000000000000000000000000000000,32'b11000000011110000000000000000000,32'b00011000000000000000000000000000,32'b00000011111000000000000000000000,32'b00000000000000000000000111000000,32'b00000000000000000000000000011111,32'b00000000000000000000011111000011,32'b00000000000000000000000000111111,32'b00000111110000110000000000000111,32'b00000111110011111101111111111111,32'b00011101100011111110000000011111,32'b01111111100011111110111000000000,32'b11100111111011111110000000000000,32'b11100011111111110111000000000000,32'b11110011110010101111100000000000,32'b11111110001111111111111000000000,32'b11000011101111010111111000000000,32'b11011000100111001101111111111100,32'b11111111100001011111111001111111,32'b11100000001000111110101111111111,32'b11100000000000000000000011110001,32'b11100000000000000000010011111110,32'b11110000000000000000000110111100,32'b11100000000000000000000000001110,32'b01100000000000000000000000011110,32'b11100000000000000000000000000100,32'b11100011111000000000000000000111,32'b10111111111111000000000000001111,32'b11011111100110111000000000011111,32'b11011111101111111000000000011000,32'b00100001100111111010000000011001,32'b00000111111111111000000000011100};
assign input_o[89] = {32'b00000000110001101100001100000000,32'b00000000010001111100000110111000,32'b00000000010000011100000001110000,32'b00000000010000010100000000111111,32'b00000000000000001100000000111110,32'b00000000100000000000000000111110,32'b00000000000000000000000000000100,32'b00000000000001111100000000000011,32'b00000000000001111100000000000111,32'b00000000000000111111000000000100,32'b00000001001111111111110000000000,32'b00000000001111001110110000011000,32'b00000000011110100000111011111110,32'b00000000011011100000101111111100,32'b00000000011110000001111111111100,32'b00000000010010000011111111111110,32'b00000100110111111000110011110000,32'b00000000111111111111110001111111,32'b00000000001111110101110001100100,32'b00000000000001111111110001111110,32'b00000000000000100111100000111010,32'b00000000000000100111100000100010,32'b00000000000000100111100000101010,32'b00000000000000100011000001101110,32'b00000001000000111011010000100011,32'b00000001000000111111100010011111,32'b00000001000000011111010000000110,32'b00000001000000000000000000000000,32'b00000001000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[90] = {32'b00000000000000000000000000000000,32'b11111111111111111111111111000000,32'b00000111000111000000000001111000,32'b11111111111111111111111101110000,32'b11111111000111110100000000000000,32'b00000000000000000000000010000010,32'b00000000000000000000000000000000,32'b10000000000000000000000000000000,32'b11110000000000000000000000000000,32'b00010000000000000000000000000000,32'b10000000000000000000000000000000,32'b00111000000000000000000000000000,32'b00000111100000000000000000000000,32'b00000000000000111000000000000000,32'b00000000001111010000000000000010,32'b00000000000011110000000000000000,32'b00000000000000011110000000000000,32'b00000000000001111100110000000100,32'b00000000000001111111111000000000,32'b00000000000001000010000100000100,32'b00000000000001111100000011101000,32'b00000000000111101111100000000011,32'b00000000000111111111110000000000,32'b00000000000110110111111100000000,32'b00000000000011111001111000000000,32'b00000000000011100000000000000000,32'b00000000000001100000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000111111000};
assign input_o[91] = {32'b00000000000000000000000000000000,32'b00000000000111000000000111111100,32'b00000000000000000001111111000010,32'b00000000000000000001110011000000,32'b00000001111000000000111111000000,32'b00000111111100000000011101000000,32'b00001110111100000000000010000000,32'b00000100111100000000111100000000,32'b00001111111100000000011100001110,32'b00001110111101000000000001100000,32'b00011110101101111000000000001000,32'b10011001000001111100000000000000,32'b00001100000000010110000000000000,32'b00001100000000000011100000001000,32'b00010110000000000001100000000000,32'b00000110001101000000100000010000,32'b00100110001100000000111111001000,32'b00000010010100000000001110000000,32'b11000010010011000000011110000000,32'b00000001101110111000000000000000,32'b10000000111111111100000000000111,32'b00000000011000000000000000000010,32'b00000000000000000000000000000001,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000011100000,32'b00000000000000000000000010100000,32'b00000000000000000000001111100000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[92] = {32'b11000000000000000000001000010000,32'b11100000000000000000010100001000,32'b11100000000000000000000000000000,32'b01010000000000000000001000000000,32'b10110000000000111000001100000000,32'b01010000000000011000001100000000,32'b00010000000000111000011110000000,32'b00000000000001110111000111000000,32'b00000000000001111011100000000000,32'b00000000000000101110111110100000,32'b00001000011000000000001100110010,32'b00000100001100111100011111100000,32'b00000000001011100100001111010000,32'b00000000001110011100000111100000,32'b00000000000111001100111111111100,32'b00000000000011001100100001011000,32'b00000000000000000110110000111100,32'b00000000000000000010010010010100,32'b00000000000000000011010010100000,32'b00000000000000000001001011100000,32'b00000000000000000001101011100000,32'b00000000000000000000111010000000,32'b00000000000000000000010101100000,32'b00000000000000000000010101100000,32'b00000000000000000000010000000000,32'b00000000000000000000111100000000,32'b00000000000000000000100010000000,32'b00000000000000000001000000000000,32'b00000000000000000001000010000000,32'b00000000000000000010000000000000,32'b00000000000000000100000000000000,32'b00000000000000000100000000000000};
assign input_o[93] = {32'b00000000000000000000000000000000,32'b00000000000000000000111111000000,32'b00000000000000000001111111100000,32'b00000000000000000000110000110000,32'b00000000000000000000110000011110,32'b00000000000000000101100000001110,32'b00000000001110001110000000001100,32'b00000000000001111111100000001000,32'b00000000001110110000000000001110,32'b00000000001111000000011110001110,32'b11111111111000000000010000001010,32'b00000000000000000000010000001100,32'b00001100000000000000000000001100,32'b00000001110000000000000000001100,32'b11111111100000111000011000101000,32'b11111100110000010000000000101111,32'b00000000000000000011111000100011,32'b11111111111110111111111111100000,32'b11111111111100000000000001110011,32'b00000000000000000000001011100100,32'b00000000000000000011100000111110,32'b00000000000000000000001000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000011,32'b00000000000000000000000000000011,32'b00000000000000000000000000000000};
assign input_o[94] = {32'b00000000000000000000000000000000,32'b01100000000000000000111110000000,32'b00010000000000000000010000000000,32'b00010000000000000000010000000000,32'b11000000000000000000000100000000,32'b11100000000000000000000000000000,32'b11110000000000000000000010000000,32'b11110000000000000000000000000000,32'b11111000000001111000000000000000,32'b11111100000011110001100000000000,32'b11111111011110111110000000000000,32'b01111100000111111111101000000000,32'b11111110001110001101101000000000,32'b11000000111100001000111000000000,32'b10000001100001110000111110000000,32'b10000001100000000001000000000000,32'b00000000000000000000111000000000,32'b00000000000000000000111000000000,32'b00000000111000000000011000000000,32'b01000001011001000000000000000000,32'b01000000001111000000000000000000,32'b00000000011111000000000000000000,32'b10000011111111111100000000000000,32'b10000000111111111100000000000000,32'b10000000111111000000000000000000,32'b00000000111011000000000000000000,32'b00000000010001000000000000000000,32'b00000000110000111000000000000000,32'b00000000110000011110000000000000,32'b00000000110000000011100000000000,32'b00000000100000000000010000000000,32'b00000000100000000000000000000000};
assign input_o[95] = {32'b00000000000000000000001100010110,32'b00000000000000000000000111111110,32'b00000000000000000000000001110010,32'b01000000000000000000000000011101,32'b00000000000000000000000000000110,32'b01000000000000111111100000000011,32'b01000000000000110011100000000000,32'b01000000000000011111000000000000,32'b10000000001111111111000000000000,32'b10000000011110011110000000000000,32'b00000000011000000110000000000000,32'b00000000011000001111000000001111,32'b00000000011000011111010000001111,32'b00000000011000001110010000001111,32'b00000000011111101111010001111110,32'b00000000011110101010011011111100,32'b00000000011111001011110001111000,32'b00000000001110111111110011111000,32'b00000000000101100111111111111000,32'b00000000001101000110001110000000,32'b00000000001101001110001110100000,32'b00000000001101001110011111111111,32'b00000000001101111100001111111011,32'b00000000001101111000000001010000,32'b00000000001111111000000000010000,32'b00000000001111111000000000011111,32'b00000000001111111110000000011111,32'b00000000000111110111110000011111,32'b00000000000001111111110000001101,32'b00000000000000000000000000001100,32'b00000000000000000000000000001111,32'b00001110000000000000000000000001};
assign input_o[96] = {32'b00000000000100101010000000000000,32'b00001100000100101010000000000000,32'b10011011000000111110010000001000,32'b11111110000000111111010000000000,32'b10001111000000111111000000000000,32'b00000000000000101010100000000000,32'b11111111100000101010100000000000,32'b00000011101110011010100000000000,32'b00111111111100011010000000000000,32'b00000000001111101010100000000000,32'b11110000000010111011000000000000,32'b00010001000011100011111111000000,32'b00001111000001100000000000111000,32'b00010011100111100110000000000000,32'b00001000000011111110000000001111,32'b00000100000011111110000011111111,32'b00000000000011111100000111110000,32'b00000000000011111000001101111111,32'b00000000000001111101111110000000,32'b00000001111101111011000000111111,32'b00000000111111111000000000000011,32'b01111110011101110011000000000000,32'b00000000000111101111100000000000,32'b00000000110000111000011111111111,32'b00000000000000011110000000000000,32'b00000000000000000111000000001111,32'b00000000000100000001111011111110,32'b11111111111100000000011111101111,32'b00000111111100111110000111111111,32'b00000000000010011111100001111110,32'b10000000000011111110111000000001,32'b11110011110000001111110000000001};
assign input_o[97] = {32'b11000000000000000000000000010000,32'b10011000000000000000000000011000,32'b11011000000000010000000000010000,32'b11000000000000010000000000001110,32'b11000000000000010000000000000111,32'b11000000000000000000000000000000,32'b11110000000000000000000000000000,32'b11111100000000000001110000000000,32'b11000110000000000000101110000000,32'b11000000110000000000000111110000,32'b11010001111000000000000111111110,32'b11000011111000000000000000110111,32'b11000000010100000000011100000000,32'b11000000001111111110011101110000,32'b11000000000001000000100000000000,32'b11000000000000000000100000000000,32'b11000000000000000000101000000000,32'b11000000000000011110011111000000,32'b11000000000000010001111111000000,32'b11000000000001001000001111000000,32'b11111111010000111111111111000000,32'b11111111111100011110011010000000,32'b11000110001100001111101000000000,32'b11110000001111100100100011000000,32'b11000000111111111111110011000000,32'b11000000000000011111110000000011,32'b11000000000000000001111000011000,32'b11000000000000000000001000000000,32'b11000000000000000000000000000000,32'b11000000000000000000000000000000,32'b11000000000000000000000000000000,32'b11000000000000000000000000000000};
assign input_o[98] = {32'b00000000100000000000000000000000,32'b00000000100000000000000000000000,32'b00000000111111111000000000000000,32'b00000000011111000000000000000000,32'b00000000000111000110000000000000,32'b00000000000011111111110000000000,32'b00000000000001110111011000000000,32'b00000000000111111011111110000000,32'b00000000000010001000011110000000,32'b00000001110011001111001110000000,32'b00000011111111000111110111100000,32'b00000001110111000111110000000000,32'b00000000011111000001110000000000,32'b00000000000100000011100000000000,32'b00000000000000000000100000000000,32'b00000000000000000000000000000000,32'b00000000000000000100000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000111000000000000,32'b00000000000000000100000000000000,32'b00000000000000110001100000000000,32'b00000000000000100010000000000000,32'b00000000000000100010000000000000,32'b00000000000000000000000000000000,32'b00000000000000000110000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
assign input_o[99] = {32'b00000000000000000001100001000010,32'b00000000000000000001111010000110,32'b00000000000000000000111000110110,32'b00000000000000000000101100011110,32'b00000000000000000001100111011011,32'b00000000000000000011111111110010,32'b00000000000000000011110011011100,32'b00000000000000000011000010111100,32'b00000000000000000111000000100000,32'b00000000000000000111000000000000,32'b00000000000000000111101111100000,32'b00000000000000000011101111100000,32'b00000000000000000011111101110000,32'b00000000000000000011000111011000,32'b00000000000000000111100111111000,32'b00000000000000111110110111111000,32'b00000000000111111110000000110000,32'b00000000011110111100000000000000,32'b00000000111101110000000000000011,32'b00000001111111000000000000011111,32'b00000001110100000000000000111110,32'b11111111111111111111111111110100,32'b11111111111111111111111110100000,32'b01111011111111111111110111100000,32'b11111111111111111111111111100100,32'b11111111111111111111111111100100,32'b11111111111111111111111011000010,32'b10111111001001111111011110000001,32'b00011110010111001100101100000000,32'b00000110011110011000011100000000,32'b00000110011111111010011011000000,32'b00000110110111010000000000000000};
endmodule
