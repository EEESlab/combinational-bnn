/* Module: parameters
 * Author: Manuele Rusci - manuele.rusci@unibo.it
 * Description: BNN net32 model weights.
 */

 module parameters
(
	output logic [15:0][0:0][8:0] weight_o_0,
	output logic [15:0][3:0] threshold_o_0,
	output logic [15:0][1:0] sign_o_0,
	output logic [31:0][15:0][8:0] weight_o_1,
	output logic [31:0][7:0] threshold_o_1,
	output logic [31:0][1:0] sign_o_1,
	output logic [47:0][31:0][8:0] weight_o_2,
	output logic [47:0][8:0] threshold_o_2,
	output logic [47:0][1:0] sign_o_2,
	output logic [63:0][47:0][8:0] weight_o_3,
	output logic [63:0][8:0] threshold_o_3,
	output logic [63:0][1:0] sign_o_3,
	output logic [63:0][255:0] weight_o_5,
	output logic [63:0][8:0] threshold_o_5,
	output logic [63:0][1:0] sign_o_5,
	output logic [3:0][63:0] weight_o_6
);
assign threshold_o_0[15:0] = {4'd4,4'd6,4'd6,4'd6,4'd5,4'd6,4'd5,4'd5,4'd6,4'd6,4'd5,4'd5,4'd6,4'd5,4'd6,4'd4};
assign sign_o_0[15:0] = {2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1};
assign weight_o_0[15:0] = {{9'b111011111},{9'b010101100},{9'b001000110},{9'b010111000},{9'b010011101},{9'b100001010},{9'b101100111},{9'b101011100},{9'b100100010},{9'b111001001},{9'b111011100},{9'b101111110},{9'b100010011},{9'b001110101},{9'b110001010},{9'b111111011}};
assign threshold_o_1[31:0] = {8'd79,8'd75,8'd78,8'd79,8'd79,8'd77,8'd79,8'd77,8'd76,8'd77,8'd79,8'd76,8'd76,8'd76,8'd75,8'd73,8'd77,8'd78,8'd79,8'd78,8'd75,8'd79,8'd78,8'd79,8'd79,8'd79,8'd74,8'd80,8'd80,8'd78,8'd77,8'd76};
assign sign_o_1[31:0] = {2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1};
assign weight_o_1[31:0] = {{9'b101001010,9'b000000001,9'b010000101,9'b010011100,9'b100000010,9'b001101010,9'b111010100,9'b101001010,9'b100001101,9'b010101000,9'b111101000,9'b011000010,9'b010101100,9'b000001000,9'b100000111,9'b100111100},{9'b111101100,9'b111000100,9'b011111111,9'b111001111,9'b010001010,9'b101010010,9'b011110100,9'b011110100,9'b101101011,9'b111101111,9'b111100001,9'b001101000,9'b111110011,9'b101101001,9'b101011000,9'b011111111},{9'b100111110,9'b011000000,9'b101010101,9'b100000010,9'b000111111,9'b010110100,9'b010011011,9'b100011000,9'b010101101,9'b111100010,9'b101011001,9'b111011110,9'b110011111,9'b101001011,9'b100100010,9'b110110101},{9'b001110111,9'b001110011,9'b011111101,9'b010001111,9'b100011100,9'b001011011,9'b000110010,9'b110000101,9'b010010011,9'b101111000,9'b110110101,9'b000010010,9'b000011110,9'b011010111,9'b000010001,9'b101110100},{9'b100011011,9'b001001001,9'b000001000,9'b100110010,9'b111011011,9'b101110100,9'b001000010,9'b111001011,9'b011100000,9'b000000001,9'b101001011,9'b100011011,9'b110011001,9'b010110011,9'b100100001,9'b010011111},{9'b111011111,9'b001000000,9'b111000000,9'b000101000,9'b011000000,9'b000100000,9'b001000110,9'b100010011,9'b001001110,9'b000010011,9'b110111101,9'b110011100,9'b001111110,9'b011100000,9'b100010111,9'b001110011},{9'b010100100,9'b110111001,9'b001101011,9'b001000000,9'b110011110,9'b110011011,9'b101010011,9'b101101111,9'b001110001,9'b001110000,9'b001010100,9'b101010110,9'b010100110,9'b110111111,9'b110000011,9'b001010101},{9'b111000110,9'b011001000,9'b111010111,9'b111001011,9'b000111100,9'b001000000,9'b110110010,9'b010010010,9'b001010001,9'b001010110,9'b000111100,9'b100110001,9'b100100111,9'b101010000,9'b000001110,9'b010111111},{9'b110111101,9'b001011111,9'b100010110,9'b110011011,9'b111111110,9'b011111011,9'b101110110,9'b111110011,9'b000000011,9'b000010000,9'b111100111,9'b001001101,9'b000100010,9'b000100101,9'b100100111,9'b111001000},{9'b111100010,9'b010010101,9'b000000010,9'b000001000,9'b101001101,9'b110010111,9'b010000100,9'b011101010,9'b000110100,9'b101011110,9'b110001001,9'b110011000,9'b101111010,9'b101000001,9'b001001110,9'b011111101},{9'b001011111,9'b000001000,9'b111111111,9'b110110011,9'b001010100,9'b111001100,9'b000111010,9'b000110110,9'b100000000,9'b101010011,9'b100101111,9'b000100011,9'b110101100,9'b111110000,9'b001000011,9'b100001111},{9'b000101100,9'b100000001,9'b001110111,9'b111011101,9'b111101110,9'b000101001,9'b001111000,9'b100000010,9'b010100000,9'b110111101,9'b110111000,9'b110001101,9'b000000000,9'b111000001,9'b100011110,9'b011000111},{9'b010110101,9'b111110111,9'b000101101,9'b010111101,9'b011111011,9'b100101101,9'b001000100,9'b101111010,9'b110110111,9'b101010111,9'b010010001,9'b000010001,9'b000100010,9'b110101111,9'b010111110,9'b011010001},{9'b010110011,9'b011011110,9'b010000110,9'b100100010,9'b110110110,9'b110001010,9'b101111001,9'b000001000,9'b101000011,9'b101101000,9'b000100001,9'b001111110,9'b011111011,9'b111111001,9'b100001110,9'b111111010},{9'b010011001,9'b110011011,9'b110110101,9'b110111111,9'b101111111,9'b001011101,9'b110110001,9'b001001011,9'b111110111,9'b010010101,9'b000101001,9'b011010001,9'b011010010,9'b000101101,9'b111111111,9'b010010101},{9'b111101101,9'b111111100,9'b100110100,9'b011011011,9'b000101001,9'b100100000,9'b010010100,9'b100011100,9'b110001011,9'b001011010,9'b011111111,9'b101000111,9'b110010111,9'b001110011,9'b010111010,9'b000111001},{9'b011010001,9'b000001011,9'b010011001,9'b100001000,9'b110011110,9'b001110010,9'b111001110,9'b001001110,9'b011111111,9'b011001000,9'b111011001,9'b101111101,9'b111110101,9'b011101101,9'b011111101,9'b111001000},{9'b000001111,9'b101100001,9'b111011100,9'b001001001,9'b000000111,9'b110110000,9'b011001001,9'b100111001,9'b000100100,9'b001010111,9'b010011110,9'b010001001,9'b101000000,9'b111101001,9'b011001111,9'b011110000},{9'b110100011,9'b111000000,9'b011111101,9'b111000110,9'b100000111,9'b000110000,9'b100011111,9'b100100001,9'b001111010,9'b011001100,9'b110001000,9'b101000001,9'b001100100,9'b101100011,9'b001010010,9'b111101001},{9'b001011010,9'b101101101,9'b101010001,9'b100000101,9'b011110010,9'b110111110,9'b111100000,9'b011000000,9'b111101110,9'b011010111,9'b101000101,9'b100111001,9'b101100011,9'b110001000,9'b101111000,9'b010001000},{9'b011110011,9'b110101111,9'b010010000,9'b000001010,9'b011010100,9'b111001110,9'b011001010,9'b000110011,9'b110011111,9'b010100110,9'b001101101,9'b011111010,9'b010111111,9'b110010000,9'b111111101,9'b100111101},{9'b110001110,9'b010101000,9'b000110110,9'b010010110,9'b000011010,9'b111011010,9'b111111100,9'b011111000,9'b000010111,9'b101001011,9'b101111110,9'b011110000,9'b010000010,9'b111111000,9'b010000000,9'b111011100},{9'b111111001,9'b000001000,9'b110110100,9'b100011011,9'b100001001,9'b101010010,9'b000101001,9'b010111001,9'b110110100,9'b111111100,9'b100111001,9'b011001000,9'b101011011,9'b011111100,9'b111000100,9'b001101000},{9'b000000011,9'b111101100,9'b110111110,9'b101010100,9'b100011011,9'b100001110,9'b000000000,9'b010101000,9'b101011111,9'b001111110,9'b110110011,9'b011001101,9'b001010001,9'b011111101,9'b010000011,9'b000010011},{9'b110100101,9'b000000101,9'b101001111,9'b100110000,9'b111010001,9'b001111101,9'b011101100,9'b000100000,9'b011111010,9'b110011011,9'b100111000,9'b010010000,9'b111011111,9'b001001101,9'b010001100,9'b111000101},{9'b100101110,9'b001101000,9'b010001001,9'b100100100,9'b010000000,9'b101011101,9'b000111100,9'b010101111,9'b011011101,9'b100100110,9'b111110110,9'b111100111,9'b101101011,9'b100101100,9'b000101000,9'b100101100},{9'b100010110,9'b111111111,9'b001000100,9'b101100111,9'b001110011,9'b011100010,9'b011001010,9'b001001101,9'b101010101,9'b100010100,9'b110111110,9'b100110010,9'b000110101,9'b011011000,9'b001110000,9'b111100100},{9'b101011010,9'b000110100,9'b111100111,9'b011001000,9'b110001100,9'b100001111,9'b101010010,9'b010001010,9'b011010111,9'b101010000,9'b001111100,9'b001000000,9'b101000111,9'b111000111,9'b100101110,9'b111000111},{9'b110110100,9'b001011000,9'b011101111,9'b001000100,9'b010110000,9'b101001011,9'b100110010,9'b000101011,9'b100001001,9'b100110111,9'b011000100,9'b000100011,9'b111100001,9'b011100011,9'b000100100,9'b010100011},{9'b110100000,9'b010111101,9'b101100110,9'b111110100,9'b011010101,9'b111111011,9'b010011111,9'b000111110,9'b011110110,9'b000100001,9'b001111010,9'b011011101,9'b011000000,9'b010000110,9'b100001111,9'b000100010},{9'b110110001,9'b110110100,9'b010001001,9'b001101011,9'b110001100,9'b011001011,9'b111010001,9'b010000010,9'b000111101,9'b011100000,9'b101100101,9'b110100101,9'b010010111,9'b000000000,9'b010010110,9'b110110101},{9'b110100001,9'b100110011,9'b010111101,9'b011011100,9'b110101000,9'b001011101,9'b000110100,9'b111100011,9'b111111010,9'b111010111,9'b011100110,9'b111101110,9'b110110110,9'b001100110,9'b111000111,9'b101000110}};
assign threshold_o_2[47:0] = {9'd152,9'd153,9'd151,9'd157,9'd151,9'd151,9'd152,9'd154,9'd159,9'd151,9'd153,9'd151,9'd150,9'd148,9'd151,9'd156,9'd155,9'd151,9'd152,9'd162,9'd154,9'd155,9'd155,9'd153,9'd152,9'd157,9'd149,9'd150,9'd152,9'd148,9'd157,9'd156,9'd157,9'd151,9'd152,9'd157,9'd152,9'd151,9'd151,9'd150,9'd156,9'd155,9'd150,9'd156,9'd149,9'd151,9'd152,9'd149};
assign sign_o_2[47:0] = {2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1};
assign weight_o_2[47:0] = {{9'b100100010,9'b100111010,9'b000111011,9'b011011001,9'b111101111,9'b001001111,9'b001111011,9'b001000101,9'b000000000,9'b101011111,9'b010110010,9'b100100000,9'b111011000,9'b101111111,9'b111111111,9'b100010000,9'b101011111,9'b001001101,9'b110100100,9'b011001010,9'b010010111,9'b001001010,9'b101000011,9'b001110001,9'b110010111,9'b010011101,9'b111011010,9'b110101110,9'b001010011,9'b000011111,9'b000001111,9'b111001011},{9'b000100100,9'b101110100,9'b010011110,9'b010011111,9'b110101010,9'b110011101,9'b000010001,9'b000010011,9'b010010101,9'b010110110,9'b010100100,9'b110111011,9'b101101101,9'b000010010,9'b110111100,9'b011100110,9'b010010001,9'b101101110,9'b110100001,9'b011111100,9'b100000001,9'b100010100,9'b111100110,9'b101101110,9'b000001010,9'b010011010,9'b010110111,9'b001001101,9'b101011111,9'b100000000,9'b011011011,9'b100010111},{9'b110001001,9'b110111111,9'b000110100,9'b010010100,9'b011010110,9'b011011110,9'b101001010,9'b101101110,9'b000011010,9'b000010001,9'b110111110,9'b111100001,9'b010000010,9'b010001111,9'b111110001,9'b101001000,9'b011100010,9'b110110101,9'b111100111,9'b100100000,9'b101001111,9'b001011010,9'b001010110,9'b101100000,9'b100101111,9'b101000011,9'b100111110,9'b110100101,9'b100101011,9'b000001100,9'b010111001,9'b000001011},{9'b001111001,9'b000010101,9'b110111011,9'b010001101,9'b110000000,9'b010010100,9'b010000101,9'b111000110,9'b010010000,9'b110111001,9'b011001001,9'b010011001,9'b010111100,9'b100011100,9'b101011100,9'b011001010,9'b001011000,9'b110010100,9'b000100011,9'b100010111,9'b010101000,9'b101001111,9'b100011000,9'b111110011,9'b100111101,9'b011000011,9'b100000001,9'b101011011,9'b001111111,9'b010100111,9'b000000100,9'b000111100},{9'b001001110,9'b100111101,9'b000100000,9'b001001100,9'b010111100,9'b001110001,9'b111000010,9'b111111011,9'b011011000,9'b000000100,9'b111101110,9'b010111111,9'b110101110,9'b100110111,9'b111000111,9'b110011000,9'b010000000,9'b110001100,9'b111011111,9'b111000011,9'b100000000,9'b010011110,9'b101111110,9'b110100011,9'b110000100,9'b100100011,9'b101111110,9'b110000011,9'b110001110,9'b110110101,9'b010010000,9'b100100101},{9'b101101011,9'b011110101,9'b111111000,9'b001001101,9'b100101111,9'b111001001,9'b110110110,9'b111100110,9'b110111100,9'b000111101,9'b110110111,9'b000101000,9'b000100001,9'b101100101,9'b000000000,9'b001111011,9'b100001100,9'b111100101,9'b101011011,9'b001100000,9'b110100110,9'b000110000,9'b000011011,9'b001001000,9'b010011011,9'b011110110,9'b110001010,9'b111010100,9'b111000101,9'b000000111,9'b010011101,9'b100110100},{9'b011001111,9'b111000011,9'b110111111,9'b000101011,9'b011110000,9'b110111101,9'b010101000,9'b000011111,9'b110000111,9'b101111011,9'b001110110,9'b001100100,9'b110000010,9'b010110100,9'b010110000,9'b101011000,9'b111100011,9'b000110000,9'b110111011,9'b010000010,9'b000011110,9'b011000110,9'b101111000,9'b110101001,9'b011110011,9'b100001011,9'b100010000,9'b011100111,9'b111011110,9'b100010011,9'b101010111,9'b111101110},{9'b111100110,9'b010011001,9'b010011010,9'b011101001,9'b010000010,9'b110110000,9'b111101011,9'b001101011,9'b110011101,9'b111110011,9'b101010000,9'b010110010,9'b110010011,9'b110010001,9'b100010110,9'b000010010,9'b100110001,9'b000110110,9'b001110000,9'b001010000,9'b010011110,9'b010110010,9'b110100110,9'b111010111,9'b101000000,9'b011011111,9'b101001101,9'b100101111,9'b101110101,9'b001000001,9'b011101100,9'b011100001},{9'b011111100,9'b010000001,9'b000000010,9'b000101110,9'b011100010,9'b000000000,9'b100110011,9'b100000100,9'b101110100,9'b011000001,9'b100000000,9'b101100101,9'b011001110,9'b010000011,9'b100110111,9'b110001101,9'b011111110,9'b110011000,9'b110110010,9'b010111011,9'b101000101,9'b011110000,9'b010011000,9'b110101110,9'b101111010,9'b000111000,9'b110011100,9'b010101000,9'b110110001,9'b011011111,9'b001100100,9'b000010010},{9'b100101010,9'b001101101,9'b110111111,9'b101011010,9'b110010100,9'b001001101,9'b110001100,9'b000000001,9'b101001000,9'b101110011,9'b100010110,9'b000010000,9'b000100010,9'b100111011,9'b111000111,9'b000001011,9'b110111111,9'b101110010,9'b010111101,9'b101100100,9'b101111111,9'b101011111,9'b001110101,9'b010110000,9'b110011100,9'b011100111,9'b100001101,9'b101010011,9'b101101111,9'b111101011,9'b100001001,9'b110101101},{9'b000001000,9'b010111101,9'b101010100,9'b010010010,9'b101100101,9'b000001110,9'b110110110,9'b010000111,9'b000101110,9'b000011001,9'b100101101,9'b011111001,9'b110000100,9'b101110010,9'b111111010,9'b001001101,9'b101110111,9'b100101011,9'b011111111,9'b101001010,9'b000100000,9'b100111100,9'b110101100,9'b111111111,9'b000111000,9'b110010110,9'b000100101,9'b100111000,9'b101110001,9'b111100011,9'b000011011,9'b111111011},{9'b101011001,9'b000010100,9'b110101001,9'b000111010,9'b101101100,9'b101110001,9'b110110101,9'b111101111,9'b010000000,9'b010001010,9'b100011000,9'b101110111,9'b100010010,9'b110100100,9'b111011100,9'b101100010,9'b100100100,9'b001101101,9'b101000001,9'b000000100,9'b000111000,9'b111110001,9'b101101111,9'b011011100,9'b000111001,9'b110010111,9'b100101000,9'b011000101,9'b110111010,9'b010110110,9'b110110111,9'b010101110},{9'b110111100,9'b011101100,9'b001010101,9'b011110000,9'b001000110,9'b001101111,9'b101001100,9'b110100101,9'b110111101,9'b001100011,9'b011011101,9'b110011011,9'b010001011,9'b100001001,9'b001011001,9'b011010110,9'b001101010,9'b110011011,9'b001110111,9'b000110000,9'b001001000,9'b111010011,9'b011011110,9'b000101010,9'b111010111,9'b110111001,9'b100100101,9'b000000110,9'b011010111,9'b000110010,9'b111100010,9'b110110001},{9'b010010000,9'b010100101,9'b100110011,9'b110111101,9'b100110111,9'b101000110,9'b111010111,9'b101111011,9'b100100001,9'b101101110,9'b000000001,9'b101101101,9'b111101000,9'b000100011,9'b001111011,9'b100111101,9'b000011001,9'b101010001,9'b010010111,9'b101101111,9'b110101110,9'b101101000,9'b100011111,9'b101101101,9'b001110111,9'b100101101,9'b111101010,9'b111001001,9'b110111011,9'b010100001,9'b110111111,9'b110111111},{9'b001011100,9'b001111010,9'b100111110,9'b101111111,9'b000111000,9'b111111111,9'b001011011,9'b110110010,9'b000000110,9'b100111100,9'b100110110,9'b010101111,9'b000001100,9'b011101110,9'b110100010,9'b011111000,9'b100111110,9'b110010100,9'b101101001,9'b000000111,9'b010010101,9'b111110011,9'b110100000,9'b000101001,9'b001101111,9'b001111111,9'b111001110,9'b100000111,9'b101011111,9'b000000011,9'b001001111,9'b000011011},{9'b110111110,9'b000010000,9'b101011101,9'b000010111,9'b110000010,9'b111100110,9'b010111001,9'b010100110,9'b111101100,9'b101110111,9'b011000010,9'b010000001,9'b110010001,9'b000001110,9'b100011100,9'b010010011,9'b000000100,9'b000001000,9'b000110010,9'b110100011,9'b000001000,9'b111011110,9'b010110010,9'b110111011,9'b110100000,9'b101000111,9'b001000110,9'b010101110,9'b100111111,9'b010000010,9'b001101100,9'b000101000},{9'b100110011,9'b011111000,9'b101011111,9'b100000010,9'b110000101,9'b100001011,9'b110101000,9'b001010011,9'b101011010,9'b001010100,9'b100100011,9'b111110000,9'b000100000,9'b111001011,9'b010000000,9'b000001000,9'b110110001,9'b000101000,9'b101010011,9'b101100110,9'b010011100,9'b000111010,9'b010000000,9'b101101100,9'b111011110,9'b100011000,9'b100000000,9'b001010101,9'b110011100,9'b111011001,9'b101111110,9'b111011101},{9'b111101101,9'b110101101,9'b110111001,9'b000110000,9'b110110000,9'b010110110,9'b101111111,9'b000111101,9'b000001000,9'b110111110,9'b000110101,9'b011000110,9'b101010101,9'b000110010,9'b100111010,9'b111110101,9'b011111100,9'b001000000,9'b100110110,9'b111000011,9'b101111101,9'b110100110,9'b110000010,9'b111100001,9'b001011111,9'b111111001,9'b101010000,9'b001011111,9'b101011100,9'b000011101,9'b110111110,9'b000101110},{9'b001010111,9'b101100000,9'b101111000,9'b110100111,9'b001110001,9'b100000011,9'b010111010,9'b010011000,9'b001100010,9'b001101110,9'b000100001,9'b101101101,9'b111111111,9'b001010000,9'b011100010,9'b100000111,9'b100110000,9'b101101011,9'b010110111,9'b111000011,9'b101010101,9'b000110001,9'b101101010,9'b001011011,9'b100110110,9'b100111111,9'b011110101,9'b000101111,9'b000000011,9'b001001010,9'b111010010,9'b110000011},{9'b011110101,9'b001000110,9'b010010010,9'b100001001,9'b111000101,9'b010000000,9'b000101110,9'b011000000,9'b111110011,9'b000000000,9'b000000000,9'b101100000,9'b111001100,9'b111001000,9'b010110011,9'b010010110,9'b110101010,9'b000000001,9'b000000001,9'b010001101,9'b010110001,9'b110010000,9'b001100100,9'b000010011,9'b001100001,9'b011000000,9'b111000010,9'b000011111,9'b001001110,9'b111111111,9'b001011000,9'b000010111},{9'b111111000,9'b100000000,9'b001000111,9'b110000000,9'b110100111,9'b100001011,9'b000001001,9'b011011101,9'b000101111,9'b111001000,9'b011110111,9'b000100011,9'b101000011,9'b001100111,9'b000101001,9'b010000111,9'b001100010,9'b100010000,9'b110110100,9'b000110000,9'b011100010,9'b011100111,9'b010100000,9'b011101101,9'b101100011,9'b010001000,9'b000010000,9'b111110101,9'b011110001,9'b110111110,9'b101010001,9'b101001110},{9'b000010101,9'b100110101,9'b111100100,9'b100101101,9'b010000000,9'b000100000,9'b011011011,9'b101011001,9'b100111100,9'b000110101,9'b110000000,9'b110111010,9'b011110010,9'b111001000,9'b010111101,9'b101000111,9'b001100010,9'b010010101,9'b100001111,9'b010011110,9'b110100001,9'b101001110,9'b100000000,9'b010000111,9'b000000111,9'b110010010,9'b100101110,9'b010000001,9'b010001001,9'b010011111,9'b000001111,9'b110101111},{9'b100101100,9'b010111010,9'b001010001,9'b010101110,9'b110111110,9'b011011001,9'b010001000,9'b010101101,9'b001010100,9'b101110011,9'b000010100,9'b101001100,9'b000010101,9'b011000001,9'b010110010,9'b001011001,9'b010011011,9'b100010011,9'b101110110,9'b100000000,9'b011011011,9'b000111100,9'b110111110,9'b110000010,9'b111110100,9'b101001101,9'b010000100,9'b111100010,9'b110101101,9'b010110111,9'b100110100,9'b010101110},{9'b111010111,9'b111000110,9'b011101101,9'b010010101,9'b011110000,9'b110100000,9'b111000000,9'b001100000,9'b111111000,9'b111111110,9'b000001001,9'b000111000,9'b100111000,9'b110011000,9'b001000111,9'b000101010,9'b000111110,9'b010001001,9'b001010001,9'b011111111,9'b101011111,9'b100010101,9'b000001101,9'b100000001,9'b101110001,9'b111111011,9'b111110110,9'b000001011,9'b001000111,9'b011001000,9'b011011011,9'b001000110},{9'b001101011,9'b110101000,9'b111101010,9'b011101011,9'b110010100,9'b011101001,9'b011110111,9'b111000010,9'b000011101,9'b110101010,9'b100000001,9'b001000000,9'b000100011,9'b110110000,9'b100111010,9'b110101000,9'b111111111,9'b011110111,9'b001000000,9'b111101111,9'b111011100,9'b110110001,9'b111110100,9'b110010001,9'b011101000,9'b111110011,9'b110110110,9'b001011000,9'b111111010,9'b111101010,9'b110110000,9'b110011001},{9'b001000101,9'b000101111,9'b011000001,9'b011101101,9'b001010101,9'b000000000,9'b000010011,9'b000000110,9'b010111001,9'b011000001,9'b000101011,9'b000100000,9'b100101000,9'b000001111,9'b111110001,9'b010111111,9'b110100010,9'b101010011,9'b101010100,9'b011010010,9'b110111111,9'b010000010,9'b011110100,9'b100110010,9'b011000000,9'b011101001,9'b000001111,9'b101000101,9'b011010010,9'b011111100,9'b010000011,9'b100111000},{9'b101111001,9'b001000001,9'b111011001,9'b010101111,9'b100101011,9'b110111111,9'b000000101,9'b101101101,9'b111100001,9'b101011111,9'b000001011,9'b111000111,9'b110001011,9'b111000101,9'b110001011,9'b100001111,9'b100001011,9'b110101100,9'b011000100,9'b100010110,9'b011001011,9'b001011011,9'b101111011,9'b011110010,9'b111111111,9'b011101001,9'b001001011,9'b100001000,9'b001110110,9'b010010000,9'b011010111,9'b001110101},{9'b000001110,9'b011111011,9'b001111101,9'b100111111,9'b111001111,9'b011101111,9'b000001001,9'b011100111,9'b100011010,9'b001101101,9'b011111011,9'b111000000,9'b010011101,9'b011001011,9'b101000110,9'b011101011,9'b011111100,9'b011001011,9'b011011011,9'b111100010,9'b001010010,9'b011001011,9'b010011000,9'b101011010,9'b111011001,9'b001111111,9'b111110110,9'b111011101,9'b111111001,9'b001101111,9'b101110111,9'b101011100},{9'b010111111,9'b101111000,9'b011111010,9'b110101000,9'b011100100,9'b101011100,9'b001101101,9'b111010001,9'b001111101,9'b001011010,9'b011010001,9'b000001000,9'b000001010,9'b001111010,9'b101100010,9'b000111101,9'b001111110,9'b010110011,9'b111101100,9'b100101010,9'b001011000,9'b000111001,9'b101010011,9'b101110011,9'b111111101,9'b011101111,9'b110000101,9'b011011011,9'b110010100,9'b011000110,9'b100110111,9'b000010000},{9'b101010101,9'b011101011,9'b101010111,9'b010110100,9'b011110010,9'b101101011,9'b111011111,9'b000111001,9'b001000011,9'b111001000,9'b101011011,9'b001001101,9'b011100001,9'b101011101,9'b101111111,9'b001011100,9'b111101011,9'b010111111,9'b111111111,9'b110100111,9'b101011111,9'b011100001,9'b011101111,9'b011110101,9'b000110111,9'b010111110,9'b001000000,9'b000111110,9'b110111011,9'b000101001,9'b111010101,9'b110001111},{9'b100011010,9'b000111111,9'b010011101,9'b011001000,9'b011010000,9'b010001000,9'b111101100,9'b111101100,9'b111010010,9'b001010010,9'b011010110,9'b101101000,9'b110000000,9'b111001010,9'b110011101,9'b011001001,9'b010001010,9'b010000000,9'b001111100,9'b100111110,9'b101000011,9'b100011001,9'b011001000,9'b110111110,9'b100001001,9'b001100000,9'b010011110,9'b110011001,9'b110100111,9'b101110111,9'b010111000,9'b010001111},{9'b110111110,9'b000100110,9'b011011101,9'b110110010,9'b000000110,9'b111111101,9'b010001000,9'b010000101,9'b111011011,9'b110011110,9'b111000111,9'b111110010,9'b111010000,9'b100000000,9'b001000000,9'b101010011,9'b101000100,9'b101000111,9'b010111010,9'b000001100,9'b000010000,9'b101000000,9'b100000010,9'b000010000,9'b000011101,9'b100100011,9'b011100111,9'b000101001,9'b000010000,9'b100000010,9'b001110011,9'b000001000},{9'b010000101,9'b101111100,9'b111010000,9'b000010001,9'b011011100,9'b001000100,9'b010100110,9'b000011010,9'b000110001,9'b100000001,9'b001000110,9'b000100001,9'b011110110,9'b110000010,9'b100111010,9'b000100010,9'b110000011,9'b001110000,9'b001010101,9'b111100100,9'b100000011,9'b101010001,9'b011100100,9'b110111011,9'b000111111,9'b110000000,9'b111001000,9'b010101001,9'b110110011,9'b000011010,9'b101010011,9'b110110101},{9'b011000001,9'b110101101,9'b011001111,9'b100011110,9'b100111000,9'b010011000,9'b101011110,9'b100101100,9'b011010000,9'b111010110,9'b000000100,9'b000001000,9'b011110000,9'b111101111,9'b011110110,9'b011001110,9'b101111010,9'b100100010,9'b001100100,9'b111110100,9'b101111111,9'b111010111,9'b001110011,9'b000110111,9'b011111010,9'b110110110,9'b000001110,9'b100001011,9'b100101010,9'b111101111,9'b010011011,9'b110000011},{9'b100110011,9'b110111011,9'b111111000,9'b100101000,9'b000000101,9'b001010011,9'b001111100,9'b010011100,9'b000010110,9'b001111001,9'b011111101,9'b111010001,9'b001000001,9'b111111110,9'b010011001,9'b000010000,9'b111101111,9'b000000000,9'b011011111,9'b010001100,9'b011111110,9'b101111011,9'b111011000,9'b011110000,9'b111110111,9'b011001100,9'b000010100,9'b111110111,9'b001111111,9'b010000011,9'b001001110,9'b001011011},{9'b111001100,9'b001001110,9'b100000100,9'b110010011,9'b000100100,9'b101100000,9'b110011000,9'b101110111,9'b011111111,9'b010000100,9'b011010000,9'b111111001,9'b000101110,9'b001101111,9'b001100001,9'b010000101,9'b010111010,9'b100101000,9'b010000000,9'b110010011,9'b000100110,9'b010100110,9'b010000000,9'b011011100,9'b001000001,9'b111110010,9'b101100101,9'b000010001,9'b011010011,9'b010110000,9'b001001001,9'b010010010},{9'b111100010,9'b110000011,9'b100111001,9'b010001101,9'b100001010,9'b001111011,9'b101010010,9'b111111111,9'b001100010,9'b011000100,9'b101110010,9'b000001011,9'b000000000,9'b011001011,9'b000001010,9'b110010000,9'b101000011,9'b011110010,9'b110111010,9'b110010010,9'b001111011,9'b110110110,9'b001100111,9'b011010100,9'b011001101,9'b100000000,9'b001000100,9'b111111111,9'b010111101,9'b111100111,9'b011111100,9'b100001011},{9'b100000011,9'b000011000,9'b111111110,9'b010101110,9'b001011000,9'b010011000,9'b111010011,9'b110111101,9'b000100110,9'b100010010,9'b001101001,9'b100100011,9'b100000001,9'b100101001,9'b011011000,9'b000001001,9'b011111000,9'b000100001,9'b100111110,9'b110100010,9'b111111101,9'b011111100,9'b001111011,9'b110101001,9'b101011001,9'b001011110,9'b100000000,9'b111111111,9'b111011110,9'b011111111,9'b100111101,9'b000111101},{9'b110110001,9'b010011101,9'b111111011,9'b000000100,9'b111111101,9'b111101110,9'b101100111,9'b011011110,9'b001000000,9'b110011101,9'b001100111,9'b010110100,9'b101000010,9'b101100110,9'b011010101,9'b001101101,9'b010011111,9'b000000110,9'b001110100,9'b000011010,9'b111111111,9'b110000011,9'b111001111,9'b001011100,9'b010101110,9'b001100111,9'b111001101,9'b011101000,9'b111100110,9'b010100000,9'b001100001,9'b000100000},{9'b100010001,9'b100010000,9'b011111010,9'b011111111,9'b110101101,9'b111111011,9'b011000010,9'b011001111,9'b001000000,9'b101111001,9'b011001100,9'b010110101,9'b000011101,9'b110001111,9'b100001111,9'b100110110,9'b011110000,9'b000001001,9'b101101001,9'b000110011,9'b101011010,9'b110011100,9'b001111000,9'b000000000,9'b011111001,9'b111101111,9'b101011110,9'b011101111,9'b111011000,9'b001100011,9'b101010100,9'b101100011},{9'b111000011,9'b100111100,9'b110100111,9'b000100001,9'b100101011,9'b010111110,9'b100111010,9'b000000000,9'b100000101,9'b000111001,9'b100000000,9'b111000100,9'b000000000,9'b000110011,9'b001111110,9'b101001001,9'b111111101,9'b000100000,9'b110000001,9'b000101011,9'b111111011,9'b100001100,9'b001010110,9'b011111001,9'b011101111,9'b001101011,9'b001010011,9'b100111001,9'b000010000,9'b100001001,9'b000001001,9'b111011011},{9'b110000011,9'b100100111,9'b000111110,9'b011000100,9'b010101100,9'b110101000,9'b010010100,9'b011111111,9'b100110111,9'b001000110,9'b111111000,9'b111111111,9'b011000110,9'b100110010,9'b101011100,9'b100010111,9'b110000110,9'b001001010,9'b001011001,9'b010000101,9'b000001001,9'b010110111,9'b000001000,9'b011000001,9'b000001110,9'b000000010,9'b101110011,9'b111001111,9'b001101000,9'b111000010,9'b111010000,9'b101001010},{9'b001001111,9'b100000000,9'b110011110,9'b001111101,9'b101011011,9'b001010011,9'b001100010,9'b101111000,9'b011011001,9'b110101111,9'b110010010,9'b010110101,9'b100111111,9'b110000000,9'b001110100,9'b100011000,9'b000000100,9'b111011111,9'b011000100,9'b100010111,9'b110101110,9'b000101111,9'b010010100,9'b000000111,9'b100000100,9'b001100010,9'b011111111,9'b000000101,9'b110101101,9'b110000011,9'b011101100,9'b101001101},{9'b000110000,9'b111110100,9'b000101001,9'b110101110,9'b000011101,9'b001000101,9'b011010000,9'b100101100,9'b010001000,9'b010010011,9'b000001001,9'b101110101,9'b111111010,9'b011000100,9'b111111111,9'b000111010,9'b010010000,9'b011010100,9'b000010111,9'b110111110,9'b001011111,9'b111110011,9'b010100110,9'b010111111,9'b100010111,9'b001110101,9'b111101100,9'b000010011,9'b000110110,9'b000010010,9'b001110000,9'b000011101},{9'b011011110,9'b111110011,9'b101110001,9'b111011111,9'b100110001,9'b010101001,9'b110011001,9'b010000100,9'b000111011,9'b101000110,9'b101010101,9'b011101111,9'b110001111,9'b111110001,9'b111111110,9'b000100110,9'b110111011,9'b101110100,9'b101101101,9'b000010010,9'b111010010,9'b011111110,9'b101110100,9'b111111110,9'b110011100,9'b100110101,9'b100110011,9'b001000000,9'b011100101,9'b100110110,9'b111000000,9'b111010100},{9'b100001100,9'b011011011,9'b011011110,9'b000101101,9'b100101100,9'b111101110,9'b101110011,9'b111101111,9'b101001101,9'b101101100,9'b011110101,9'b000111110,9'b111101100,9'b010011001,9'b000101010,9'b101001111,9'b101011101,9'b011000010,9'b100000000,9'b010000001,9'b000010100,9'b011010001,9'b101110000,9'b011101000,9'b000001001,9'b110100101,9'b000010001,9'b110110011,9'b000110000,9'b011100110,9'b100000101,9'b000000001},{9'b111010111,9'b001000000,9'b001101111,9'b000100101,9'b001111011,9'b100011111,9'b110110010,9'b110110111,9'b100100110,9'b011101101,9'b000000011,9'b101100100,9'b110000100,9'b011111010,9'b001000010,9'b111111000,9'b011000101,9'b011011111,9'b100011010,9'b111011101,9'b110100011,9'b001000010,9'b110101010,9'b011111110,9'b000011111,9'b010100111,9'b100001000,9'b000100000,9'b110111111,9'b010010011,9'b100100110,9'b000010101},{9'b000010111,9'b001111110,9'b011111111,9'b101110100,9'b010100111,9'b100111111,9'b110110111,9'b110110111,9'b100000110,9'b101010110,9'b100110111,9'b111011110,9'b110110010,9'b100101101,9'b101111010,9'b101000101,9'b110111100,9'b100011100,9'b111111111,9'b000000110,9'b000100100,9'b110100110,9'b010011011,9'b011100101,9'b010000111,9'b011101100,9'b001100100,9'b111101111,9'b101110110,9'b100111110,9'b110100111,9'b111101110}};
assign threshold_o_3[63:0] = {9'd228,9'd218,9'd234,9'd227,9'd226,9'd222,9'd227,9'd232,9'd227,9'd225,9'd233,9'd225,9'd243,9'd227,9'd226,9'd223,9'd225,9'd235,9'd219,9'd221,9'd236,9'd232,9'd226,9'd225,9'd234,9'd231,9'd233,9'd236,9'd222,9'd236,9'd233,9'd227,9'd227,9'd241,9'd238,9'd234,9'd237,9'd228,9'd232,9'd244,9'd230,9'd220,9'd240,9'd230,9'd229,9'd241,9'd232,9'd227,9'd233,9'd232,9'd243,9'd223,9'd237,9'd227,9'd231,9'd222,9'd225,9'd233,9'd226,9'd242,9'd236,9'd235,9'd249,9'd242};
assign sign_o_3[63:0] = {2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1};
assign weight_o_3[63:0] = {{9'b001001100,9'b001001110,9'b010001011,9'b111111001,9'b111001110,9'b101001011,9'b101000011,9'b001000110,9'b011011001,9'b011010001,9'b000011000,9'b111101001,9'b011111101,9'b000010101,9'b011101011,9'b000000101,9'b111111001,9'b010100000,9'b100100000,9'b110101100,9'b110111011,9'b001000111,9'b001010100,9'b001001010,9'b001100000,9'b000011100,9'b001110101,9'b100110001,9'b000110111,9'b001111000,9'b101100101,9'b101011101,9'b100111001,9'b001001011,9'b000011011,9'b001110010,9'b011111111,9'b000011000,9'b011100100,9'b110001101,9'b101101111,9'b111011011,9'b001001110,9'b000011011,9'b101111110,9'b011001010,9'b110100001,9'b100111011},{9'b010101001,9'b101011101,9'b111111111,9'b000101000,9'b110010111,9'b010110000,9'b111111011,9'b100100111,9'b101111101,9'b101101101,9'b001100110,9'b101011110,9'b101101110,9'b100010100,9'b110011011,9'b011100111,9'b110101100,9'b001111101,9'b110100100,9'b100011001,9'b101001001,9'b010010000,9'b101111111,9'b001111111,9'b111011110,9'b010011001,9'b100111110,9'b110101101,9'b110101111,9'b101100111,9'b101010010,9'b011001011,9'b100110100,9'b010111110,9'b001110101,9'b000010011,9'b110101111,9'b010001111,9'b101100101,9'b111011101,9'b100111000,9'b011010011,9'b111001110,9'b101101111,9'b101110111,9'b001011111,9'b010000001,9'b100010000},{9'b000100100,9'b100101010,9'b011011101,9'b111111001,9'b001011111,9'b100000010,9'b100110111,9'b111001000,9'b010111001,9'b011010010,9'b000011111,9'b100110010,9'b010100001,9'b101110110,9'b001100011,9'b100010000,9'b110010010,9'b001011101,9'b100111101,9'b000011100,9'b110010101,9'b100111100,9'b001110011,9'b111101100,9'b010001001,9'b001001010,9'b011101111,9'b011110101,9'b001000001,9'b000010011,9'b010110010,9'b000101111,9'b100111100,9'b000011011,9'b000011000,9'b001111110,9'b100110000,9'b000000011,9'b010101111,9'b001101110,9'b101010001,9'b101101000,9'b011101100,9'b000011010,9'b001110100,9'b111110010,9'b100110001,9'b000111010},{9'b000110001,9'b001101001,9'b111011011,9'b100010100,9'b110011001,9'b110110000,9'b111010010,9'b001001111,9'b100100010,9'b110001011,9'b101001011,9'b101111011,9'b011011111,9'b000000110,9'b010101111,9'b011100111,9'b000111110,9'b011101110,9'b101101000,9'b000110001,9'b110101111,9'b111101011,9'b001001011,9'b100011101,9'b101001000,9'b110010001,9'b011001010,9'b110010000,9'b101110110,9'b101011000,9'b110010011,9'b101101100,9'b010101101,9'b001101000,9'b110110010,9'b011011101,9'b111111111,9'b110110010,9'b010000010,9'b101001101,9'b000000000,9'b100111000,9'b011101101,9'b010001001,9'b001011000,9'b011001011,9'b010101111,9'b000111000},{9'b011100101,9'b010100110,9'b111111001,9'b110011011,9'b111010011,9'b110010011,9'b001001011,9'b001111110,9'b111111011,9'b000000100,9'b000111010,9'b010010010,9'b100111001,9'b111000010,9'b111110110,9'b111111000,9'b010010111,9'b101001111,9'b101011011,9'b101000010,9'b101111011,9'b110100011,9'b010110100,9'b110000111,9'b000010000,9'b010100010,9'b110101001,9'b000111111,9'b000010101,9'b010110111,9'b010000101,9'b111111001,9'b110001001,9'b000001010,9'b111001100,9'b101110010,9'b101000000,9'b000011000,9'b000111000,9'b110001110,9'b000011111,9'b011101111,9'b111101011,9'b100100101,9'b011011110,9'b011111101,9'b111010000,9'b011001110},{9'b101100110,9'b111110111,9'b110000101,9'b101011010,9'b001001101,9'b111001000,9'b111100000,9'b101101010,9'b000011101,9'b111001111,9'b010010000,9'b100100010,9'b101001110,9'b011111011,9'b011100101,9'b000000101,9'b000000111,9'b101100001,9'b100110010,9'b001000011,9'b001101010,9'b010001110,9'b111011001,9'b110011011,9'b111110011,9'b001110010,9'b101000111,9'b001011001,9'b101101000,9'b101011101,9'b100111011,9'b111000011,9'b011010001,9'b111011101,9'b111101001,9'b001011010,9'b111100001,9'b111011100,9'b101000111,9'b101001001,9'b111101001,9'b111011011,9'b111000110,9'b110011111,9'b111101000,9'b111110100,9'b110000111,9'b011010010},{9'b010000010,9'b001101101,9'b111111001,9'b011000011,9'b010101011,9'b011100010,9'b100001011,9'b101101100,9'b010010010,9'b110111110,9'b111010100,9'b110010110,9'b011011011,9'b110101010,9'b011101100,9'b010000011,9'b110110011,9'b011110001,9'b010010000,9'b010010010,9'b111001111,9'b000000011,9'b111111111,9'b010110000,9'b111110100,9'b000001010,9'b011011110,9'b011011011,9'b011011011,9'b011001110,9'b110001110,9'b011000010,9'b110010010,9'b001111110,9'b111101011,9'b100100110,9'b111000001,9'b011010110,9'b111001111,9'b111111110,9'b100110001,9'b101101011,9'b101110111,9'b010110111,9'b011101111,9'b110101001,9'b000010010,9'b111010110},{9'b011001110,9'b000010001,9'b010010100,9'b011111110,9'b101100111,9'b110111101,9'b001100101,9'b111111001,9'b001101111,9'b010010000,9'b011011000,9'b000110000,9'b110111001,9'b111101000,9'b010011010,9'b000100111,9'b001100100,9'b000000001,9'b000111011,9'b100000111,9'b101100110,9'b111011111,9'b000000001,9'b001100011,9'b000000110,9'b001111100,9'b001100101,9'b101011010,9'b000110101,9'b001101010,9'b001111010,9'b000101111,9'b001011010,9'b011100100,9'b000010011,9'b110110000,9'b000100101,9'b100000000,9'b110010001,9'b100111010,9'b110101111,9'b011111110,9'b100011001,9'b001000001,9'b000111001,9'b110111110,9'b101001000,9'b011010011},{9'b000111001,9'b110011101,9'b110111111,9'b010001100,9'b110010010,9'b110001011,9'b111000111,9'b110111010,9'b111111001,9'b011110110,9'b001001011,9'b010101101,9'b111110100,9'b111000110,9'b110000111,9'b000000001,9'b110000001,9'b111100001,9'b010011001,9'b011000011,9'b010111000,9'b111001001,9'b001010010,9'b110100000,9'b100101011,9'b111111100,9'b000110110,9'b111010010,9'b001011110,9'b000000110,9'b111001010,9'b110111101,9'b110010010,9'b011011011,9'b110101010,9'b001001101,9'b011010001,9'b100100101,9'b001100010,9'b100111101,9'b000101011,9'b100101101,9'b111111001,9'b000101111,9'b101011110,9'b000111010,9'b110010000,9'b100010011},{9'b001100100,9'b100111110,9'b111101010,9'b010101010,9'b110010110,9'b100010000,9'b100110011,9'b000100110,9'b000010011,9'b101110011,9'b100110110,9'b011101110,9'b001011001,9'b100110110,9'b100111001,9'b110010001,9'b111101000,9'b011010000,9'b110000100,9'b110010001,9'b000011011,9'b001000110,9'b101101110,9'b111011010,9'b110001110,9'b100010110,9'b111101010,9'b101010010,9'b011011011,9'b001000100,9'b011111111,9'b001011001,9'b001000010,9'b100111100,9'b011010111,9'b111110111,9'b011011011,9'b011011011,9'b101010111,9'b111101011,9'b001011110,9'b010110010,9'b100101011,9'b100110100,9'b010111111,9'b101010110,9'b001011101,9'b000010110},{9'b110101100,9'b000011010,9'b110100110,9'b101101000,9'b110000000,9'b000000010,9'b000100101,9'b001000100,9'b101110100,9'b100111011,9'b000110011,9'b011110111,9'b000100010,9'b001111100,9'b001111011,9'b111011000,9'b001111011,9'b001111000,9'b001001000,9'b100011100,9'b001010011,9'b111110000,9'b100100111,9'b111101000,9'b000001010,9'b001001011,9'b111111111,9'b100001010,9'b101001111,9'b100100011,9'b010110001,9'b100101100,9'b101011001,9'b110111001,9'b000101001,9'b100110000,9'b100111011,9'b000111010,9'b001000011,9'b100100101,9'b111111000,9'b111000001,9'b011000110,9'b110011000,9'b000101000,9'b111000000,9'b111110111,9'b100101100},{9'b110111000,9'b010100001,9'b101110010,9'b001101101,9'b110100000,9'b011011010,9'b010001110,9'b111010100,9'b010000010,9'b000111110,9'b001101111,9'b010011110,9'b111101010,9'b000011111,9'b110101111,9'b000101011,9'b100010111,9'b111111101,9'b010001100,9'b000110100,9'b110011011,9'b011010011,9'b001101111,9'b000010111,9'b111110100,9'b000000110,9'b001001111,9'b010001011,9'b001001110,9'b011101101,9'b011001110,9'b010000001,9'b000011110,9'b011111010,9'b011101111,9'b011110100,9'b000011110,9'b010000111,9'b101101111,9'b111000111,9'b110111011,9'b110110011,9'b000111101,9'b001111110,9'b001000000,9'b000111001,9'b011111110,9'b101101110},{9'b100011100,9'b010111100,9'b101010000,9'b100011101,9'b100010010,9'b011100101,9'b001110011,9'b100010000,9'b000110011,9'b001110000,9'b010000001,9'b100000000,9'b111110001,9'b000000100,9'b011110010,9'b110111011,9'b110000110,9'b001000000,9'b110010101,9'b101001111,9'b000100010,9'b001001100,9'b110010010,9'b000011100,9'b010111101,9'b001000110,9'b100100100,9'b001110110,9'b101101111,9'b011110011,9'b100000010,9'b101001011,9'b100010011,9'b000001000,9'b001110011,9'b010110100,9'b010110010,9'b000000010,9'b101100010,9'b000001010,9'b000111000,9'b011011001,9'b101110100,9'b100110000,9'b100100010,9'b011110001,9'b010111100,9'b101000000},{9'b110001001,9'b100101101,9'b000000100,9'b110111111,9'b111111100,9'b000001000,9'b000100111,9'b100101110,9'b100110010,9'b000000001,9'b110111111,9'b110011110,9'b110110111,9'b110000101,9'b010001101,9'b010101100,9'b100101010,9'b100000011,9'b010010111,9'b111011011,9'b100110110,9'b101011111,9'b101010001,9'b000001100,9'b111000000,9'b000101000,9'b011001000,9'b000100101,9'b011000101,9'b101101100,9'b100001101,9'b110110100,9'b110011011,9'b000001001,9'b101100001,9'b010001110,9'b110001011,9'b000001000,9'b001000000,9'b001010101,9'b100001010,9'b111100111,9'b101010101,9'b001110010,9'b010100010,9'b010101000,9'b010010010,9'b111100011},{9'b100110100,9'b100000101,9'b001110010,9'b110011010,9'b000000101,9'b110110010,9'b100111110,9'b110001100,9'b001110110,9'b010111010,9'b110111110,9'b110111110,9'b101100011,9'b010101101,9'b111111101,9'b011000001,9'b010000010,9'b100111111,9'b101100101,9'b011001011,9'b010101010,9'b100001111,9'b000111100,9'b111101000,9'b100110101,9'b100001111,9'b100100100,9'b110100001,9'b001111010,9'b001110101,9'b010011001,9'b001010011,9'b001001000,9'b111110000,9'b110010000,9'b100000010,9'b110010000,9'b010110011,9'b101101111,9'b101111101,9'b101011110,9'b100001011,9'b000100110,9'b011000101,9'b100100010,9'b001010000,9'b111000101,9'b110110111},{9'b101010001,9'b011000001,9'b100000011,9'b011110111,9'b101101101,9'b001001111,9'b101101111,9'b001011011,9'b011001011,9'b000100101,9'b101111000,9'b000001101,9'b101010001,9'b011001011,9'b000000001,9'b011111111,9'b010001010,9'b001101000,9'b110011011,9'b100110110,9'b100101011,9'b000111111,9'b000010111,9'b000111001,9'b000101111,9'b101011011,9'b011100111,9'b110110011,9'b001000011,9'b100001100,9'b100000000,9'b101111111,9'b101101001,9'b001000101,9'b110010111,9'b011001111,9'b011000011,9'b100000100,9'b110010001,9'b101001101,9'b111111111,9'b101101100,9'b100001011,9'b111100001,9'b111010100,9'b010000110,9'b001011111,9'b101001100},{9'b111110110,9'b000000111,9'b111110101,9'b111100101,9'b001000000,9'b101111011,9'b111001000,9'b110001111,9'b000011011,9'b101111101,9'b101010111,9'b110110000,9'b010000001,9'b011101110,9'b101111010,9'b101100101,9'b011010011,9'b011101010,9'b011000111,9'b100000110,9'b010110000,9'b000000110,9'b000111100,9'b011010011,9'b011111000,9'b000111001,9'b001111101,9'b101101001,9'b101011000,9'b101011011,9'b001011000,9'b100011000,9'b100010001,9'b111111101,9'b111001110,9'b010110110,9'b001101000,9'b101011001,9'b111011101,9'b011011010,9'b111111101,9'b010010001,9'b101100110,9'b010010110,9'b001100001,9'b100010110,9'b111110100,9'b101001000},{9'b101111011,9'b100011001,9'b100011110,9'b111101000,9'b000000110,9'b101011111,9'b110111011,9'b001001000,9'b000000101,9'b010011010,9'b000101101,9'b111111111,9'b010101000,9'b010111000,9'b011111000,9'b001001000,9'b100010011,9'b110111011,9'b010000000,9'b010101011,9'b001000001,9'b101011001,9'b000001000,9'b111000010,9'b011111010,9'b011100111,9'b001000010,9'b000000000,9'b100011010,9'b000101011,9'b010111011,9'b111001000,9'b000000000,9'b001001011,9'b011111011,9'b110101000,9'b111000010,9'b111010011,9'b110011011,9'b000111000,9'b100001011,9'b000000100,9'b100110111,9'b001101101,9'b011001111,9'b111011110,9'b000111001,9'b100000101},{9'b000101010,9'b011011010,9'b011110110,9'b111101111,9'b011111110,9'b000101100,9'b000100011,9'b100000010,9'b010101110,9'b010011111,9'b001111110,9'b111111111,9'b111110111,9'b011101010,9'b001111111,9'b111100000,9'b110101010,9'b011101010,9'b110000111,9'b111111101,9'b100011011,9'b110111001,9'b010010101,9'b110011001,9'b011000111,9'b110101101,9'b011010100,9'b110101101,9'b001111101,9'b101111111,9'b111000000,9'b100000001,9'b101000011,9'b001011111,9'b100100110,9'b110110010,9'b001100111,9'b111110101,9'b010000101,9'b100000111,9'b000000110,9'b110100101,9'b111111001,9'b010110001,9'b100101010,9'b011001111,9'b111100011,9'b110100010},{9'b101110010,9'b111100110,9'b111111011,9'b111011011,9'b111000011,9'b011000011,9'b011101000,9'b111101101,9'b010101011,9'b111010100,9'b001001001,9'b010110010,9'b111110011,9'b100101011,9'b111110110,9'b000000111,9'b000011011,9'b111100111,9'b110111010,9'b000000011,9'b101100010,9'b010010001,9'b111111011,9'b110100101,9'b110111000,9'b100010000,9'b111101001,9'b011100001,9'b111011110,9'b110110010,9'b101010000,9'b000110001,9'b000010010,9'b100000110,9'b111111100,9'b010111010,9'b110001011,9'b011010000,9'b100110011,9'b111011010,9'b101000010,9'b101011011,9'b101010101,9'b101110110,9'b111001101,9'b101001111,9'b111010110,9'b110101011},{9'b011110010,9'b000000101,9'b110111001,9'b011001110,9'b110000000,9'b111111110,9'b110100100,9'b011001111,9'b100100110,9'b110010111,9'b001001010,9'b011000100,9'b100010110,9'b100101000,9'b000110000,9'b001010110,9'b100110000,9'b111011000,9'b000010000,9'b111110100,9'b111011001,9'b010001001,9'b000001010,9'b001100100,9'b011111100,9'b100110101,9'b011001000,9'b000100000,9'b010101111,9'b001110110,9'b100100010,9'b101110000,9'b011001000,9'b010011001,9'b010110000,9'b100100101,9'b111101110,9'b010011110,9'b110101101,9'b001100100,9'b000001001,9'b111110001,9'b011001001,9'b001011010,9'b000011011,9'b010101011,9'b111101000,9'b100100000},{9'b000010000,9'b000001001,9'b111111001,9'b010010110,9'b101011010,9'b101010000,9'b011001001,9'b011101001,9'b101100110,9'b000111011,9'b010000000,9'b011001101,9'b000011010,9'b001110001,9'b111000101,9'b100010111,9'b010110101,9'b010111011,9'b011101100,9'b110110111,9'b001010111,9'b110111011,9'b011001001,9'b100111101,9'b000101101,9'b000010001,9'b101101001,9'b000010000,9'b000100100,9'b001011000,9'b101010010,9'b001110010,9'b011110100,9'b010011011,9'b011111011,9'b011100100,9'b001110110,9'b011110010,9'b111010100,9'b011001111,9'b101111000,9'b111011010,9'b110001101,9'b010101001,9'b011110000,9'b010100000,9'b101010110,9'b011000001},{9'b110000010,9'b011011111,9'b110111011,9'b010011000,9'b100101100,9'b000000100,9'b100001110,9'b001100000,9'b010001111,9'b011111110,9'b000110100,9'b010110110,9'b110001011,9'b010000110,9'b000011100,9'b001100000,9'b111110110,9'b001001100,9'b001001101,9'b111111100,9'b101001010,9'b111011101,9'b110010110,9'b000111110,9'b000000101,9'b100011010,9'b111011111,9'b111100111,9'b110001111,9'b000011011,9'b010010010,9'b111010011,9'b001110100,9'b000110111,9'b011101011,9'b001101010,9'b111010110,9'b000101100,9'b100001001,9'b100101000,9'b110110110,9'b111000011,9'b101100010,9'b010111110,9'b111100000,9'b111000010,9'b100111000,9'b101000101},{9'b011101010,9'b111001111,9'b111111111,9'b000111000,9'b110110011,9'b110111101,9'b110000101,9'b101011011,9'b010101001,9'b100011111,9'b010111010,9'b110101110,9'b110011100,9'b100111011,9'b111101111,9'b010101100,9'b111011100,9'b100101101,9'b011100101,9'b011100001,9'b110110010,9'b100110100,9'b111010110,9'b010110101,9'b110000001,9'b010011100,9'b000010111,9'b010011101,9'b100010110,9'b001011000,9'b100010111,9'b110011000,9'b101010100,9'b100000101,9'b111101001,9'b100101001,9'b000010010,9'b000001110,9'b001000111,9'b111110111,9'b000000110,9'b111100001,9'b100010010,9'b010000000,9'b100110011,9'b100001011,9'b000110100,9'b111001001},{9'b010010010,9'b100001101,9'b100010010,9'b011000001,9'b010010110,9'b000010101,9'b111010011,9'b100101011,9'b010110001,9'b100111100,9'b100100001,9'b000010110,9'b001000010,9'b100100110,9'b110101001,9'b001001011,9'b011011011,9'b001100000,9'b011101010,9'b111110000,9'b101010011,9'b111111110,9'b100100010,9'b111110000,9'b100111011,9'b100011100,9'b100100100,9'b010100001,9'b110001111,9'b100001110,9'b010011110,9'b001001101,9'b011011001,9'b110110011,9'b001100110,9'b111100110,9'b010011010,9'b011011010,9'b001011000,9'b001000101,9'b000111110,9'b100000010,9'b001111000,9'b000100110,9'b110100100,9'b100000100,9'b000001101,9'b111000101},{9'b001001100,9'b001100001,9'b100111111,9'b001100000,9'b011000011,9'b000001101,9'b001001111,9'b101000001,9'b101101010,9'b101011110,9'b001110100,9'b001000100,9'b000001000,9'b011111000,9'b010100001,9'b000011101,9'b011111000,9'b110101101,9'b001100110,9'b001011000,9'b001011110,9'b101010001,9'b111010000,9'b011101111,9'b000011110,9'b101001011,9'b101011111,9'b011011011,9'b101001011,9'b000111111,9'b001100010,9'b110011001,9'b001100100,9'b101010001,9'b001010111,9'b001010101,9'b010011001,9'b001100111,9'b001001001,9'b111000001,9'b111110010,9'b111001001,9'b011000010,9'b001110010,9'b101100101,9'b010011011,9'b000100110,9'b001100101},{9'b011011001,9'b000000101,9'b111111110,9'b001000001,9'b010000101,9'b001111000,9'b100111110,9'b101100001,9'b111100101,9'b000011011,9'b011001001,9'b001000100,9'b101110000,9'b011000100,9'b010001001,9'b011011101,9'b010100100,9'b010011010,9'b010000000,9'b110110110,9'b001111011,9'b110101000,9'b000011011,9'b110110111,9'b011011011,9'b000100111,9'b000100010,9'b001100100,9'b000110001,9'b101011011,9'b000000110,9'b101001101,9'b111011111,9'b000010111,9'b001110100,9'b111000000,9'b100011110,9'b000111110,9'b101101110,9'b110000101,9'b001100010,9'b100000000,9'b010011001,9'b000111010,9'b100100000,9'b100000100,9'b111110101,9'b110010000},{9'b111111110,9'b000100011,9'b001000010,9'b110111100,9'b010011101,9'b011001011,9'b111110001,9'b101101010,9'b100010000,9'b101100111,9'b100010010,9'b010110101,9'b000001101,9'b000000110,9'b000110001,9'b101110001,9'b111100000,9'b000101010,9'b010000111,9'b001111100,9'b000100010,9'b000000010,9'b100101000,9'b101100110,9'b000110111,9'b100100100,9'b101001111,9'b101000000,9'b100001100,9'b100101011,9'b000001000,9'b110110010,9'b110101010,9'b100000101,9'b101011100,9'b010100000,9'b000111000,9'b000011100,9'b111110100,9'b111111011,9'b110101100,9'b010000000,9'b100011110,9'b100100010,9'b011100011,9'b111101100,9'b110111010,9'b010001001},{9'b101001010,9'b110101111,9'b111000010,9'b100111111,9'b110011010,9'b110000001,9'b011011100,9'b111111101,9'b111101000,9'b111100010,9'b001101001,9'b011001100,9'b111001010,9'b110111101,9'b111000011,9'b110110110,9'b001001011,9'b111001101,9'b101110101,9'b000011000,9'b011010101,9'b110011001,9'b111010001,9'b110111000,9'b010000001,9'b000011010,9'b101010011,9'b111000101,9'b001100000,9'b011110101,9'b111111000,9'b011101100,9'b110101100,9'b110000111,9'b101100010,9'b111110111,9'b011000101,9'b111000000,9'b110000111,9'b110100101,9'b101011000,9'b011011001,9'b001111111,9'b111110010,9'b111011100,9'b101111011,9'b011101100,9'b010000000},{9'b110001000,9'b111100100,9'b110010000,9'b001000001,9'b111001111,9'b001011011,9'b011100010,9'b101101100,9'b001001010,9'b011111010,9'b011011100,9'b010000101,9'b101001110,9'b111101000,9'b011000001,9'b000001110,9'b001010111,9'b011111111,9'b001101000,9'b010011001,9'b000011111,9'b000011111,9'b000100110,9'b000100010,9'b011011100,9'b011010110,9'b100100000,9'b010000010,9'b000101101,9'b000000110,9'b000110011,9'b000100111,9'b010111011,9'b110000100,9'b010110100,9'b011100010,9'b000011110,9'b011000000,9'b101100001,9'b000000111,9'b111101100,9'b011000000,9'b110100100,9'b100110100,9'b010110110,9'b110100011,9'b001001111,9'b011110000},{9'b000111001,9'b000001000,9'b101111111,9'b111111110,9'b000000000,9'b100010010,9'b010111011,9'b001000111,9'b001100001,9'b011011010,9'b000110000,9'b001010010,9'b101000011,9'b000111100,9'b010111100,9'b101001011,9'b011111010,9'b110110100,9'b000011101,9'b111011011,9'b101101111,9'b011110010,9'b000111001,9'b011101001,9'b000011000,9'b010111001,9'b011011011,9'b010101101,9'b000111110,9'b100111010,9'b111111010,9'b000000000,9'b011000000,9'b101111000,9'b100111100,9'b101111101,9'b111111000,9'b101111010,9'b100111101,9'b100110010,9'b101101000,9'b000000101,9'b101000010,9'b001000000,9'b000011000,9'b010001001,9'b111110001,9'b100110110},{9'b011001101,9'b011000111,9'b110001001,9'b100010110,9'b001010110,9'b110110001,9'b011011011,9'b110101001,9'b011100010,9'b111110000,9'b010010000,9'b011100100,9'b100100101,9'b000101111,9'b101000001,9'b011100110,9'b000100000,9'b011011001,9'b010110100,9'b001010101,9'b011011000,9'b000001111,9'b000100010,9'b000100101,9'b110100100,9'b100110111,9'b111101111,9'b101011010,9'b111101010,9'b111111110,9'b000001010,9'b001010111,9'b001100000,9'b100110000,9'b100101100,9'b000000011,9'b101000110,9'b111010101,9'b010101111,9'b101101000,9'b101110111,9'b110000011,9'b110000101,9'b110100110,9'b010111111,9'b110100110,9'b101000111,9'b111010011},{9'b000011011,9'b011101111,9'b100100110,9'b111101000,9'b101001101,9'b011110100,9'b110110001,9'b000111011,9'b101111001,9'b001110100,9'b001001011,9'b110001001,9'b101100110,9'b010111111,9'b011011001,9'b111111000,9'b000100110,9'b100010001,9'b110011001,9'b101110100,9'b100111010,9'b000001001,9'b001000000,9'b001100101,9'b101111101,9'b100111010,9'b101000011,9'b100001000,9'b011100001,9'b001111010,9'b110101100,9'b100001101,9'b101111001,9'b100111111,9'b110001100,9'b101001101,9'b111111100,9'b110001000,9'b001100011,9'b111011111,9'b001011101,9'b011111101,9'b010000100,9'b001000010,9'b001011011,9'b010000111,9'b111110011,9'b100111000},{9'b010011101,9'b101010010,9'b100111101,9'b110101100,9'b101101100,9'b101000010,9'b000010111,9'b000000001,9'b111101000,9'b010010100,9'b111011011,9'b001000010,9'b011101000,9'b111101110,9'b111000100,9'b101000100,9'b101010000,9'b000001010,9'b010000000,9'b111101011,9'b110011000,9'b101100010,9'b000100100,9'b011000100,9'b110100000,9'b000011010,9'b100100100,9'b000110101,9'b101100110,9'b000101110,9'b110010011,9'b000010110,9'b000110100,9'b001111010,9'b100000011,9'b010111000,9'b101000100,9'b010000000,9'b001001111,9'b101001000,9'b100111110,9'b000001000,9'b011000100,9'b010001100,9'b100111000,9'b000000001,9'b101100100,9'b000001011},{9'b110010110,9'b000000111,9'b100100011,9'b000001000,9'b011100011,9'b001100111,9'b110100111,9'b010001011,9'b000111001,9'b001000000,9'b110000011,9'b011011000,9'b100110001,9'b010010010,9'b010000011,9'b001100001,9'b100101100,9'b001001000,9'b010010101,9'b010111001,9'b101100100,9'b010110010,9'b000000100,9'b000000101,9'b010000001,9'b101001111,9'b101111001,9'b000000101,9'b000100100,9'b000101000,9'b001001011,9'b110111001,9'b010010001,9'b011001011,9'b101100110,9'b010000111,9'b111010010,9'b100001100,9'b100001101,9'b100100110,9'b110101111,9'b000100011,9'b101010011,9'b010001011,9'b001000100,9'b100100110,9'b001010111,9'b011000001},{9'b011000000,9'b011100001,9'b001011000,9'b111000101,9'b110000110,9'b110001100,9'b010010100,9'b100000010,9'b100000011,9'b100001010,9'b101110110,9'b111100010,9'b010010000,9'b100100111,9'b101010010,9'b001101100,9'b111100010,9'b011001101,9'b000100100,9'b011010011,9'b010100001,9'b010100011,9'b010110100,9'b110000011,9'b101000011,9'b110010010,9'b101000000,9'b111000000,9'b011001110,9'b101000111,9'b100010111,9'b110100100,9'b000010011,9'b100010011,9'b010000001,9'b000011010,9'b111011111,9'b001101111,9'b011010010,9'b011001111,9'b001001011,9'b100000100,9'b110000101,9'b110000100,9'b111110010,9'b000000011,9'b001000111,9'b100000110},{9'b010111011,9'b001001000,9'b001010011,9'b110110010,9'b010000100,9'b110010010,9'b010110111,9'b000000011,9'b110101000,9'b010001011,9'b000000110,9'b000111110,9'b100000000,9'b000011000,9'b111111010,9'b101100000,9'b011110100,9'b101011101,9'b101001000,9'b011111100,9'b011000111,9'b001000000,9'b001001001,9'b000111010,9'b110000110,9'b011010101,9'b101110001,9'b000010010,9'b011100010,9'b000010100,9'b111010000,9'b110010100,9'b100011010,9'b011111111,9'b010010001,9'b011001000,9'b110010111,9'b001110111,9'b100001011,9'b001000000,9'b110111101,9'b001110000,9'b101001100,9'b001001000,9'b000010001,9'b111111100,9'b111101100,9'b010110011},{9'b000100110,9'b010100111,9'b001101110,9'b101111010,9'b111111001,9'b101000011,9'b001111110,9'b100011111,9'b111101000,9'b000100000,9'b010110010,9'b001001100,9'b011011011,9'b010000000,9'b100101111,9'b110011111,9'b100100001,9'b001000101,9'b110000110,9'b111101101,9'b111111000,9'b001001001,9'b011110001,9'b010000010,9'b000000011,9'b001111000,9'b110001111,9'b101001110,9'b101100011,9'b001100100,9'b110001110,9'b110101111,9'b110000100,9'b010010000,9'b000100101,9'b100000000,9'b010000000,9'b000000001,9'b101000000,9'b100001001,9'b101001101,9'b001001011,9'b111000111,9'b110010110,9'b011001111,9'b010000101,9'b110111101,9'b001000001},{9'b100000000,9'b100100100,9'b010100001,9'b111000110,9'b101001111,9'b101000101,9'b010001000,9'b000000010,9'b111110100,9'b110110010,9'b111001001,9'b010000010,9'b100101101,9'b100001001,9'b010000000,9'b110101110,9'b110000100,9'b000100000,9'b011000111,9'b011110100,9'b011100000,9'b010110001,9'b110110100,9'b010111111,9'b110000011,9'b001011100,9'b010100011,9'b100110111,9'b111011011,9'b111011011,9'b111110111,9'b001000101,9'b010110100,9'b100000000,9'b001001011,9'b110011001,9'b011001100,9'b100001000,9'b100000101,9'b100001001,9'b100000010,9'b011101010,9'b101001011,9'b101110000,9'b010110010,9'b111111010,9'b100100110,9'b001001001},{9'b010110111,9'b100010101,9'b111110010,9'b100001000,9'b011101001,9'b010000001,9'b001110000,9'b001010000,9'b010011100,9'b010011000,9'b000111111,9'b111100000,9'b011001110,9'b011110101,9'b101100000,9'b111001001,9'b110010000,9'b011111100,9'b011000111,9'b110110000,9'b011011000,9'b100010000,9'b000111000,9'b010000001,9'b001010110,9'b010111010,9'b001000000,9'b000010110,9'b010001000,9'b011110110,9'b001010000,9'b010100001,9'b000110001,9'b011111111,9'b001111000,9'b000001101,9'b001100000,9'b000011000,9'b000111001,9'b101101101,9'b100110010,9'b010000001,9'b101000011,9'b101110110,9'b001011110,9'b100000010,9'b110100001,9'b001011001},{9'b100110000,9'b101110111,9'b001110001,9'b100110010,9'b101000100,9'b100000110,9'b100111110,9'b010001100,9'b110010100,9'b111111110,9'b001110011,9'b111010111,9'b110110010,9'b000110001,9'b000101100,9'b000011010,9'b000000001,9'b000110110,9'b011110010,9'b010000000,9'b011101011,9'b010000100,9'b111111111,9'b111000100,9'b110010110,9'b100000000,9'b101111001,9'b010110100,9'b010011100,9'b001101101,9'b000110011,9'b000110000,9'b010000010,9'b011000111,9'b111111011,9'b010011111,9'b001111010,9'b110110011,9'b011011101,9'b110101101,9'b001011101,9'b101100101,9'b010010101,9'b010011010,9'b111011111,9'b111101011,9'b100110010,9'b100100110},{9'b101111001,9'b100010100,9'b101000010,9'b000111011,9'b000110000,9'b111000010,9'b111011000,9'b011101010,9'b000101110,9'b111101111,9'b011000100,9'b101111111,9'b111101100,9'b111111100,9'b110001010,9'b011100110,9'b001010001,9'b111101000,9'b111011100,9'b000111111,9'b110011101,9'b001000101,9'b111100100,9'b100100111,9'b111111101,9'b000101100,9'b110110110,9'b101110100,9'b110101001,9'b101100100,9'b001101000,9'b010000101,9'b101101101,9'b111100011,9'b111111000,9'b010010111,9'b011100111,9'b101101111,9'b111110110,9'b101101001,9'b111111111,9'b010011010,9'b100010110,9'b100110111,9'b100100000,9'b111001101,9'b111111101,9'b010100010},{9'b000010001,9'b011101011,9'b101001110,9'b111011001,9'b111111100,9'b001000110,9'b001000101,9'b001010000,9'b111111101,9'b100001100,9'b001000011,9'b011000001,9'b101000101,9'b100101011,9'b100000111,9'b000011000,9'b010000001,9'b000001101,9'b011000011,9'b011011000,9'b110111000,9'b010001011,9'b011000100,9'b010001110,9'b000000010,9'b101111110,9'b011000000,9'b001010000,9'b011001010,9'b010100000,9'b110101000,9'b011110101,9'b100001000,9'b000000001,9'b001001000,9'b011110101,9'b100000010,9'b110100001,9'b010000110,9'b100000110,9'b011100001,9'b000110111,9'b111011010,9'b111100000,9'b011110111,9'b000000000,9'b001000000,9'b001111110},{9'b000000101,9'b100100110,9'b100110111,9'b011001000,9'b101101101,9'b100000110,9'b011000010,9'b000000100,9'b111101101,9'b100111101,9'b100000000,9'b011110110,9'b110100100,9'b110000101,9'b100000010,9'b001101000,9'b111011101,9'b001001010,9'b001000100,9'b110011111,9'b100111000,9'b011011010,9'b011100010,9'b111000100,9'b010000100,9'b000111101,9'b010101010,9'b100000101,9'b111010100,9'b011000000,9'b010111110,9'b111111111,9'b101010000,9'b000100100,9'b110001110,9'b101110100,9'b011010011,9'b101000010,9'b101001101,9'b101001001,9'b000101000,9'b000010111,9'b011100100,9'b101101101,9'b000011110,9'b101010011,9'b011000000,9'b000001110},{9'b010001101,9'b111111101,9'b011100001,9'b100101010,9'b110010010,9'b010000011,9'b111110100,9'b001111001,9'b000001111,9'b100000000,9'b011010000,9'b101001100,9'b101111011,9'b000000010,9'b011101100,9'b000011111,9'b010111010,9'b011011011,9'b011110111,9'b000010111,9'b100100110,9'b101011000,9'b110011011,9'b000101110,9'b110110100,9'b010111000,9'b110001011,9'b000010010,9'b000111001,9'b101110000,9'b110100000,9'b101111110,9'b110011111,9'b110001010,9'b101100110,9'b000110011,9'b001001110,9'b001001000,9'b001000111,9'b001000110,9'b000001000,9'b100011011,9'b111011001,9'b100010111,9'b001001000,9'b101110111,9'b000101101,9'b000111010},{9'b011101101,9'b000000011,9'b011101111,9'b000101100,9'b010000011,9'b011000011,9'b000000001,9'b000001010,9'b100100001,9'b100110000,9'b001010100,9'b010010101,9'b001101101,9'b101000001,9'b000010010,9'b110011010,9'b011000011,9'b001000000,9'b001110011,9'b110111110,9'b111100110,9'b000000000,9'b001000001,9'b000010000,9'b011011000,9'b110111100,9'b010001000,9'b001000010,9'b000011001,9'b111000010,9'b111110100,9'b110000111,9'b010111110,9'b010001111,9'b010001011,9'b010011000,9'b101100110,9'b111100100,9'b110100100,9'b000100000,9'b110101010,9'b100011001,9'b101000110,9'b110010000,9'b010011010,9'b010101001,9'b100100011,9'b001011010},{9'b101110001,9'b111101000,9'b010111011,9'b001110111,9'b100010110,9'b011000001,9'b000011010,9'b001100001,9'b001110100,9'b110110010,9'b010011010,9'b110000110,9'b000001101,9'b111000110,9'b100000001,9'b100100110,9'b110100000,9'b100011011,9'b101100100,9'b101101110,9'b000010000,9'b011010010,9'b000100101,9'b110100000,9'b000100000,9'b110011101,9'b100100111,9'b010100111,9'b100010111,9'b010101010,9'b010000111,9'b011111111,9'b011110100,9'b110010100,9'b001110111,9'b110000000,9'b011001100,9'b011010110,9'b111100101,9'b010010010,9'b101110111,9'b100011010,9'b110100000,9'b100100110,9'b111100000,9'b101001111,9'b011100100,9'b011010001},{9'b100011101,9'b100100101,9'b110111110,9'b001000010,9'b111100001,9'b011000010,9'b000001001,9'b000000101,9'b111101000,9'b100111010,9'b011011110,9'b000000000,9'b001100101,9'b110010100,9'b010100101,9'b101100001,9'b101000101,9'b001010001,9'b001000110,9'b111110010,9'b100001110,9'b101110000,9'b101100100,9'b011110100,9'b001000111,9'b110111111,9'b100001101,9'b001010110,9'b101100011,9'b101100111,9'b011101000,9'b011001111,9'b000010010,9'b110110111,9'b011011111,9'b111010111,9'b101000110,9'b011100010,9'b111000010,9'b110011101,9'b001111111,9'b001000101,9'b101100000,9'b011100100,9'b001111111,9'b000100001,9'b000001000,9'b011010101},{9'b111001011,9'b100011101,9'b011100000,9'b100110011,9'b100000101,9'b110100001,9'b010110111,9'b011111001,9'b010000001,9'b110000011,9'b000111001,9'b110111101,9'b001100001,9'b010101001,9'b000011000,9'b110011010,9'b010110101,9'b010111010,9'b000010001,9'b100000011,9'b010100001,9'b000000011,9'b010011001,9'b111000001,9'b000110001,9'b000010100,9'b111111001,9'b010110011,9'b111110001,9'b011011001,9'b010011011,9'b000010011,9'b010000101,9'b010100000,9'b010111001,9'b100101010,9'b111011010,9'b011111101,9'b010111111,9'b111111011,9'b000101011,9'b110001010,9'b110100100,9'b000100001,9'b000111001,9'b001010101,9'b111101011,9'b000111011},{9'b110011111,9'b100110010,9'b011001110,9'b101111000,9'b000001010,9'b010000011,9'b010010000,9'b110110010,9'b111111000,9'b000110111,9'b101011101,9'b110100010,9'b000001011,9'b000001010,9'b110000010,9'b010010110,9'b111101100,9'b010000010,9'b010000101,9'b111001100,9'b110000100,9'b000110000,9'b111101011,9'b011101110,9'b101110001,9'b001111011,9'b110101110,9'b110010111,9'b101110110,9'b010010011,9'b110110110,9'b010000010,9'b110111000,9'b100111011,9'b011010010,9'b011110001,9'b111001100,9'b110110110,9'b110011111,9'b110010001,9'b010110010,9'b110100100,9'b100100001,9'b110111110,9'b111110000,9'b110010010,9'b100001100,9'b010000101},{9'b000111110,9'b000101111,9'b000101000,9'b110111100,9'b001000000,9'b000000110,9'b000011110,9'b001011000,9'b110010010,9'b001010100,9'b010110010,9'b000001110,9'b110001100,9'b000101100,9'b101101010,9'b100000001,9'b000000010,9'b000011010,9'b101110110,9'b101010100,9'b011111001,9'b000000000,9'b010110111,9'b100010000,9'b101110110,9'b010100110,9'b011001000,9'b000100010,9'b101110010,9'b001111000,9'b110111111,9'b101000100,9'b000111000,9'b111110110,9'b000111010,9'b001000011,9'b010011011,9'b010011110,9'b011010110,9'b000011011,9'b101111110,9'b001010000,9'b111000010,9'b111011110,9'b010100110,9'b010001010,9'b100010110,9'b000011111},{9'b010110110,9'b001111011,9'b001001010,9'b110011010,9'b111010001,9'b101100010,9'b001000100,9'b011010011,9'b101100010,9'b011100111,9'b011000111,9'b101110111,9'b110000010,9'b001101011,9'b001110111,9'b000010010,9'b001100111,9'b111111110,9'b110010011,9'b101010101,9'b000100100,9'b001111010,9'b011010110,9'b010101000,9'b111111110,9'b001000111,9'b011100101,9'b011011110,9'b011000100,9'b000110010,9'b110011111,9'b001100000,9'b001100000,9'b011111111,9'b110010111,9'b101100100,9'b101111111,9'b101110111,9'b110110001,9'b111001111,9'b011111110,9'b110101111,9'b110011001,9'b100111011,9'b011100010,9'b000111000,9'b001110110,9'b111110111},{9'b000000001,9'b110100101,9'b110001000,9'b001110101,9'b011100111,9'b100001110,9'b111000111,9'b010010100,9'b100111011,9'b000001101,9'b110001001,9'b010110101,9'b110010101,9'b100101001,9'b010001101,9'b000100111,9'b110101101,9'b110000000,9'b100110001,9'b001011001,9'b000110010,9'b000110001,9'b100001100,9'b000110100,9'b110111010,9'b000011001,9'b001001011,9'b000001110,9'b100100100,9'b000000000,9'b111110110,9'b110110101,9'b111101011,9'b001000001,9'b101000001,9'b010111010,9'b001010000,9'b110000110,9'b100000100,9'b100100001,9'b001011000,9'b010011110,9'b010001001,9'b000010001,9'b100010010,9'b110101010,9'b010111011,9'b110001111},{9'b100010000,9'b111101001,9'b011001001,9'b010011110,9'b110011010,9'b010000111,9'b000101111,9'b100001110,9'b110010000,9'b110111111,9'b110111101,9'b101111110,9'b111010110,9'b100111101,9'b111101011,9'b100100110,9'b010111010,9'b001000111,9'b000110110,9'b110101100,9'b101100101,9'b110111000,9'b111001000,9'b011001000,9'b100000111,9'b011111001,9'b101100001,9'b000010011,9'b110010001,9'b000011010,9'b010110111,9'b100101001,9'b010101100,9'b111001101,9'b010010111,9'b111110010,9'b110010011,9'b010111010,9'b111000010,9'b010000000,9'b100101000,9'b101000010,9'b011100100,9'b000111001,9'b010011001,9'b111010011,9'b000000110,9'b010100110},{9'b101101111,9'b111001010,9'b100101001,9'b111100100,9'b000110111,9'b110110101,9'b001111001,9'b010011101,9'b111011000,9'b011111011,9'b111010001,9'b000000000,9'b010000010,9'b010001011,9'b110110101,9'b111001000,9'b001000100,9'b100100010,9'b011010010,9'b011100110,9'b111000000,9'b110111111,9'b110010001,9'b000110110,9'b100110011,9'b000110010,9'b011010110,9'b111011111,9'b010001000,9'b011011010,9'b110011000,9'b100000111,9'b111000011,9'b000110011,9'b101011000,9'b000010111,9'b000111000,9'b110110010,9'b011100001,9'b110101111,9'b000011111,9'b010111101,9'b101000011,9'b011010110,9'b001001101,9'b011011101,9'b001001000,9'b101001010},{9'b011110010,9'b110000000,9'b100000110,9'b111111101,9'b100000101,9'b100101101,9'b110111000,9'b010111010,9'b000001110,9'b110010110,9'b111111001,9'b011011001,9'b011010110,9'b110010011,9'b111111011,9'b110111001,9'b101000101,9'b110100100,9'b100001010,9'b010100111,9'b111110110,9'b011111101,9'b001011010,9'b000000101,9'b011011001,9'b100110110,9'b110100111,9'b100100110,9'b101011101,9'b011101000,9'b100100100,9'b101110111,9'b001111101,9'b011011111,9'b100100000,9'b001101111,9'b111100111,9'b001100100,9'b001010110,9'b111100000,9'b010111010,9'b101101101,9'b111110011,9'b001000011,9'b010101101,9'b011111110,9'b110011111,9'b111110101},{9'b110100101,9'b101100100,9'b011110011,9'b111111100,9'b010111111,9'b001011011,9'b111000011,9'b011011111,9'b000111011,9'b010111001,9'b110110000,9'b000100000,9'b000110101,9'b111001001,9'b011111010,9'b110000100,9'b100110011,9'b011101010,9'b111011111,9'b001000001,9'b011001001,9'b001011100,9'b100111101,9'b101001110,9'b101000100,9'b000100101,9'b100101101,9'b110100011,9'b100000100,9'b110101101,9'b111100001,9'b110111101,9'b100001010,9'b100010000,9'b110010110,9'b101010010,9'b000011100,9'b110001011,9'b101010111,9'b111000101,9'b111111111,9'b111100010,9'b111000110,9'b000011000,9'b111111110,9'b000111100,9'b101100100,9'b001011010},{9'b000100000,9'b101101111,9'b001100101,9'b111000000,9'b000110010,9'b011100111,9'b101000010,9'b111100110,9'b110101000,9'b011101011,9'b010111110,9'b100000010,9'b010101111,9'b001111100,9'b010001001,9'b111110000,9'b100111001,9'b001101000,9'b100000000,9'b101011000,9'b011111000,9'b011111010,9'b111100101,9'b011100000,9'b000011010,9'b111110111,9'b101000111,9'b110000111,9'b010000000,9'b000001000,9'b111011100,9'b100000110,9'b101111000,9'b010011000,9'b010101101,9'b011011000,9'b111100000,9'b101000101,9'b101001010,9'b111000110,9'b001001100,9'b010000011,9'b001110101,9'b010001000,9'b001111110,9'b000000011,9'b110001010,9'b010110110},{9'b100010111,9'b101100001,9'b111110111,9'b100110000,9'b011001000,9'b011000110,9'b000000010,9'b100100000,9'b111101001,9'b000000110,9'b110010101,9'b001111110,9'b110000000,9'b101100011,9'b011001100,9'b111011011,9'b011011111,9'b001100110,9'b111111110,9'b001011110,9'b110000001,9'b000111100,9'b100111111,9'b101000111,9'b000001100,9'b010000001,9'b100011010,9'b100110000,9'b101011011,9'b101111111,9'b001011000,9'b000100000,9'b110110110,9'b110111011,9'b110110110,9'b011110100,9'b000011010,9'b110011101,9'b111111110,9'b101110010,9'b111111111,9'b011010110,9'b101101000,9'b100110100,9'b100110010,9'b111100100,9'b000111011,9'b010000000},{9'b101111110,9'b000011010,9'b010000010,9'b111110011,9'b000000010,9'b000101010,9'b011000010,9'b001111010,9'b100010101,9'b101110001,9'b100111010,9'b001101010,9'b001100000,9'b010100011,9'b001001110,9'b100000000,9'b101010101,9'b000000011,9'b100011011,9'b010010111,9'b101110000,9'b010010010,9'b101000101,9'b000000011,9'b100011000,9'b011010111,9'b101001101,9'b100001011,9'b010100001,9'b110111000,9'b111111010,9'b000100110,9'b010110000,9'b000001000,9'b101000010,9'b000010000,9'b100001101,9'b110110000,9'b001010111,9'b010011010,9'b011111101,9'b010010010,9'b011000001,9'b100010001,9'b010001000,9'b110100100,9'b100010101,9'b010110111},{9'b111000000,9'b101101110,9'b011001010,9'b011010101,9'b000111001,9'b110110000,9'b101000001,9'b101100110,9'b011011011,9'b110000011,9'b110111001,9'b110011100,9'b001010100,9'b101101101,9'b100110111,9'b000100100,9'b100100001,9'b000101000,9'b000111100,9'b010111101,9'b010010111,9'b111110001,9'b001000101,9'b001111110,9'b111101000,9'b100010000,9'b010001011,9'b101001111,9'b000100001,9'b000100000,9'b000001001,9'b100111000,9'b010011000,9'b011100001,9'b010000010,9'b100110100,9'b000001001,9'b110000000,9'b000000011,9'b001000000,9'b001110001,9'b101111111,9'b111110000,9'b000011011,9'b001100000,9'b111110010,9'b000001110,9'b111001100},{9'b000011000,9'b100110100,9'b001111101,9'b100011010,9'b011001101,9'b100001011,9'b001110101,9'b001001111,9'b101000100,9'b110010100,9'b111100010,9'b001001111,9'b010100001,9'b100101011,9'b001011100,9'b100110000,9'b000011001,9'b000011000,9'b110101100,9'b100000000,9'b100000010,9'b001001100,9'b110010111,9'b101101101,9'b111111111,9'b001000110,9'b000100101,9'b001110010,9'b000110100,9'b100111100,9'b010000000,9'b000011011,9'b000111000,9'b110110101,9'b001111011,9'b101100101,9'b010011001,9'b100110111,9'b111101101,9'b001111000,9'b101101011,9'b001001010,9'b111110010,9'b000111000,9'b011110011,9'b000010001,9'b100111110,9'b111101000},{9'b010101100,9'b110100000,9'b000100110,9'b110110011,9'b000100001,9'b100000100,9'b000111010,9'b100101111,9'b111010000,9'b010111100,9'b000101000,9'b011111101,9'b000100011,9'b001111100,9'b000111010,9'b111110000,9'b110100001,9'b001011100,9'b000111000,9'b011001000,9'b100010011,9'b010000000,9'b010110110,9'b001010000,9'b010011100,9'b100100101,9'b000110100,9'b000011000,9'b010111110,9'b000110011,9'b110110010,9'b010101001,9'b101110000,9'b101100101,9'b010011000,9'b000000000,9'b110010010,9'b110111010,9'b011010111,9'b000001111,9'b000011100,9'b001010100,9'b000100100,9'b001010010,9'b100100111,9'b000001100,9'b100101100,9'b000010000},{9'b001001100,9'b100100100,9'b111011101,9'b110100100,9'b101000010,9'b100011000,9'b001000010,9'b011000110,9'b100111000,9'b010010011,9'b000001010,9'b000010001,9'b001111011,9'b111100000,9'b011001000,9'b110010101,9'b100100100,9'b011101000,9'b001100110,9'b010110000,9'b000011101,9'b100111100,9'b001000100,9'b111011110,9'b000000100,9'b010110110,9'b011000100,9'b000000001,9'b101100100,9'b011001111,9'b110110100,9'b010111011,9'b000010100,9'b001000010,9'b110001100,9'b110101000,9'b000000101,9'b110100000,9'b001000110,9'b010000101,9'b100010111,9'b111011010,9'b011010100,9'b101110100,9'b001000010,9'b000101011,9'b000000100,9'b101100001}};
assign threshold_o_5[63:0] = {9'd128,9'd129,9'd125,9'd129,9'd130,9'd130,9'd129,9'd132,9'd133,9'd126,9'd129,9'd124,9'd135,9'd136,9'd130,9'd129,9'd129,9'd126,9'd129,9'd134,9'd124,9'd133,9'd124,9'd125,9'd126,9'd131,9'd123,9'd130,9'd125,9'd124,9'd129,9'd125,9'd124,9'd132,9'd130,9'd127,9'd136,9'd131,9'd127,9'd131,9'd126,9'd125,9'd126,9'd131,9'd132,9'd129,9'd135,9'd132,9'd128,9'd128,9'd131,9'd130,9'd130,9'd134,9'd131,9'd128,9'd126,9'd132,9'd129,9'd130,9'd131,9'd129,9'd127,9'd133};
assign sign_o_5[63:0] = {2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1};
assign weight_o_5[63:0] = {{1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0},{1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0},{1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0},{1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0},{1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0},{1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0},{1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0},{1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0},{1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0},{1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0},{1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1},{1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1},{1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0},{1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0},{1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1},{1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0},{1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0},{1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1},{1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1},{1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0},{1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1},{1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1},{1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0},{1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0},{1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0},{1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1},{1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0},{1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0},{1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1},{1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1},{1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1},{1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1},{1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0},{1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1},{1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1},{1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1},{1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0},{1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0},{1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1},{1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0},{1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1},{1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1},{1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0},{1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1},{1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0},{1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0},{1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0},{1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0},{1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1},{1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1},{1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1},{1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1},{1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0},{1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0},{1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1},{1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0},{1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1},{1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1},{1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1},{1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1},{1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0},{1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1},{1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1},{1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}};
assign weight_o_6[3:0] = {{1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1},{1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1},{1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1},{1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b0,1'b1}};
endmodule
